`timescale 1ns / 1ps

`include "s15850_scan.v"

module tb_s15850;
    integer fptr;
    localparam Size = 720896;
    reg [87:0] test_data [720895:0];
    integer i = 0;

    reg CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
            g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
            g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
            g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
            g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
            g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
            g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
            test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
            test_si10;

    wire g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
            g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
            g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
            g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
            g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
            g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
            g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
            g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
            g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
            g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
            g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
            g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
            g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
            g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
            g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
            g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
            test_so6, test_so7, test_so8, test_so9, test_so10;

    `define in_data {g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,           g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84, g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892, g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9, test_si10}

    s15850 inst_s15850 (
    .CK (CK),
    .g100 (g100),
    .g101 (g101),
    .g102 (g102),
    .g103 (g103),
    .g10377 (g10377),
    .g10379 (g10379),
    .g104 (g104),
    .g10455 (g10455),
    .g10457 (g10457),
    .g10459 (g10459),
    .g10461 (g10461),
    .g10463 (g10463),
    .g10465 (g10465),
    .g10628 (g10628),
    .g10801 (g10801),
    .g109 (g109),
    .g11163 (g11163),
    .g11206 (g11206),
    .g11489 (g11489),
    .g1170 (g1170),
    .g1173 (g1173),
    .g1176 (g1176),
    .g1179 (g1179),
    .g1182 (g1182),
    .g1185 (g1185),
    .g1188 (g1188),
    .g1191 (g1191),
    .g1194 (g1194),
    .g1197 (g1197),
    .g1200 (g1200),
    .g1203 (g1203),
    .g1696 (g1696),
    .g1700 (g1700),
    .g1712 (g1712),
    .g18 (g18),
    .g1957 (g1957),
    .g1960 (g1960),
    .g1961 (g1961),
    .g23 (g23),
    .g2355 (g2355),
    .g2601 (g2601),
    .g2602 (g2602),
    .g2603 (g2603),
    .g2604 (g2604),
    .g2605 (g2605),
    .g2606 (g2606),
    .g2607 (g2607),
    .g2608 (g2608),
    .g2609 (g2609),
    .g2610 (g2610),
    .g2611 (g2611),
    .g2612 (g2612),
    .g2648 (g2648),
    .g27 (g27),
    .g28 (g28),
    .g29 (g29),
    .g2986 (g2986),
    .g30 (g30),
    .g3007 (g3007),
    .g3069 (g3069),
    .g31 (g31),
    .g3327 (g3327),
    .g41 (g41),
    .g4171 (g4171),
    .g4172 (g4172),
    .g4173 (g4173),
    .g4174 (g4174),
    .g4175 (g4175),
    .g4176 (g4176),
    .g4177 (g4177),
    .g4178 (g4178),
    .g4179 (g4179),
    .g4180 (g4180),
    .g4181 (g4181),
    .g4191 (g4191),
    .g4192 (g4192),
    .g4193 (g4193),
    .g4194 (g4194),
    .g4195 (g4195),
    .g4196 (g4196),
    .g4197 (g4197),
    .g4198 (g4198),
    .g4199 (g4199),
    .g42 (g42),
    .g4200 (g4200),
    .g4201 (g4201),
    .g4202 (g4202),
    .g4203 (g4203),
    .g4204 (g4204),
    .g4205 (g4205),
    .g4206 (g4206),
    .g4207 (g4207),
    .g4208 (g4208),
    .g4209 (g4209),
    .g4210 (g4210),
    .g4211 (g4211),
    .g4212 (g4212),
    .g4213 (g4213),
    .g4214 (g4214),
    .g4215 (g4215),
    .g4216 (g4216),
    .g43 (g43),
    .g44 (g44),
    .g45 (g45),
    .g46 (g46),
    .g47 (g47),
    .g48 (g48),
    .g4887 (g4887),
    .g4888 (g4888),
    .g5101 (g5101),
    .g5105 (g5105),
    .g5658 (g5658),
    .g5659 (g5659),
    .g5816 (g5816),
    .g6253 (g6253),
    .g6254 (g6254),
    .g6255 (g6255),
    .g6256 (g6256),
    .g6257 (g6257),
    .g6258 (g6258),
    .g6259 (g6259),
    .g6260 (g6260),
    .g6261 (g6261),
    .g6262 (g6262),
    .g6263 (g6263),
    .g6264 (g6264),
    .g6265 (g6265),
    .g6266 (g6266),
    .g6267 (g6267),
    .g6268 (g6268),
    .g6269 (g6269),
    .g6270 (g6270),
    .g6271 (g6271),
    .g6272 (g6272),
    .g6273 (g6273),
    .g6274 (g6274),
    .g6275 (g6275),
    .g6276 (g6276),
    .g6277 (g6277),
    .g6278 (g6278),
    .g6279 (g6279),
    .g6280 (g6280),
    .g6281 (g6281),
    .g6282 (g6282),
    .g6283 (g6283),
    .g6284 (g6284),
    .g6285 (g6285),
    .g6842 (g6842),
    .g6920 (g6920),
    .g6926 (g6926),
    .g6932 (g6932),
    .g6942 (g6942),
    .g6949 (g6949),
    .g6955 (g6955),
    .g741 (g741),
    .g742 (g742),
    .g743 (g743),
    .g744 (g744),
    .g750 (g750),
    .g7744 (g7744),
    .g8061 (g8061),
    .g8062 (g8062),
    .g82 (g82),
    .g8271 (g8271),
    .g83 (g83),
    .g8313 (g8313),
    .g8316 (g8316),
    .g8318 (g8318),
    .g8323 (g8323),
    .g8328 (g8328),
    .g8331 (g8331),
    .g8335 (g8335),
    .g8340 (g8340),
    .g8347 (g8347),
    .g8349 (g8349),
    .g8352 (g8352),
    .g84 (g84),
    .g85 (g85),
    .g8561 (g8561),
    .g8562 (g8562),
    .g8563 (g8563),
    .g8564 (g8564),
    .g8565 (g8565),
    .g8566 (g8566),
    .g86 (g86),
    .g87 (g87),
    .g872 (g872),
    .g873 (g873),
    .g877 (g877),
    .g88 (g88),
    .g881 (g881),
    .g886 (g886),
    .g889 (g889),
    .g89 (g89),
    .g892 (g892),
    .g895 (g895),
    .g8976 (g8976),
    .g8977 (g8977),
    .g8978 (g8978),
    .g8979 (g8979),
    .g898 (g898),
    .g8980 (g8980),
    .g8981 (g8981),
    .g8982 (g8982),
    .g8983 (g8983),
    .g8984 (g8984),
    .g8985 (g8985),
    .g8986 (g8986),
    .g90 (g90),
    .g901 (g901),
    .g904 (g904),
    .g907 (g907),
    .g91 (g91),
    .g910 (g910),
    .g913 (g913),
    .g916 (g916),
    .g919 (g919),
    .g92 (g92),
    .g922 (g922),
    .g925 (g925),
    .g93 (g93),
    .g94 (g94),
    .g9451 (g9451),
    .g95 (g95),
    .g96 (g96),
    .g99 (g99),
    .g9961 (g9961),
    .test_se (test_se),
    .test_si1 (test_si1),
    .test_so1 (test_so1),
    .test_si2 (test_si2),
    .test_so2 (test_so2),
    .test_si3 (test_si3),
    .test_so3 (test_so3),
    .test_si4 (test_si4),
    .test_so4 (test_so4),
    .test_si5 (test_si5),
    .test_so5 (test_so5),
    .test_si6 (test_si6),
    .test_so6 (test_so6),
    .test_si7 (test_si7),
    .test_so7 (test_so7),
    .test_si8 (test_si8),
    .test_so8 (test_so8),
    .test_si9 (test_si9),
    .test_so9 (test_so9),
    .test_si10 (test_si10),
    .test_so10 (test_so10)
    );

    initial begin
        // $dumpfile("s15850.vcd");
        // $dumpvars(0, tb_s15850);
        fptr = $fopen("data_out.txt", "w");

        $readmemb("s15808_12samples.vec", test_data);
        for (i=0; i<Size; i = i + 1) begin
            `in_data = test_data[i]; #10;

            $fwrite(fptr, "%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d\n", inst_s15850.g100, inst_s15850.g101, inst_s15850.g102, inst_s15850.g103, inst_s15850.g104, inst_s15850.g109, inst_s15850.g1170, inst_s15850.g1173, inst_s15850.g1176, inst_s15850.g1179, inst_s15850.g1182, inst_s15850.g1185, inst_s15850.g1188, inst_s15850.g1191, inst_s15850.g1194, inst_s15850.g1197, inst_s15850.g1200, inst_s15850.g1203, inst_s15850.g1696, inst_s15850.g1700, inst_s15850.g1712, inst_s15850.g18, inst_s15850.g1960, inst_s15850.g1961, inst_s15850.g23, inst_s15850.g27, inst_s15850.g28, inst_s15850.g29, inst_s15850.g30, inst_s15850.g31, inst_s15850.g41, inst_s15850.g42, inst_s15850.g43, inst_s15850.g44, inst_s15850.g45, inst_s15850.g46, inst_s15850.g47, inst_s15850.g48, inst_s15850.g741, inst_s15850.g742, inst_s15850.g743, inst_s15850.g744, inst_s15850.g750, inst_s15850.g82, inst_s15850.g83, inst_s15850.g84, inst_s15850.g85, inst_s15850.g86, inst_s15850.g87, inst_s15850.g872, inst_s15850.g873, inst_s15850.g877, inst_s15850.g88, inst_s15850.g881, inst_s15850.g886, inst_s15850.g889, inst_s15850.g89, inst_s15850.g892, inst_s15850.g895, inst_s15850.g898, inst_s15850.g90, inst_s15850.g901, inst_s15850.g904, inst_s15850.g907, inst_s15850.g91, inst_s15850.g910, inst_s15850.g913, inst_s15850.g916, inst_s15850.g919, inst_s15850.g92, inst_s15850.g922, inst_s15850.g925, inst_s15850.g93, inst_s15850.g94, inst_s15850.g95, inst_s15850.g96, inst_s15850.g99, inst_s15850.test_se, inst_s15850.test_si1, inst_s15850.test_si2, inst_s15850.test_si3, inst_s15850.test_si4, inst_s15850.test_si5, inst_s15850.test_si6, inst_s15850.test_si7, inst_s15850.test_si8, inst_s15850.test_si9, inst_s15850.test_si10, inst_s15850.g10377, inst_s15850.g10379, inst_s15850.g10455, inst_s15850.g10457, inst_s15850.g10459, inst_s15850.g10461, inst_s15850.g10463, inst_s15850.g10465, inst_s15850.g10628, inst_s15850.g10801, inst_s15850.g11163, inst_s15850.g11206, inst_s15850.g11489, inst_s15850.g1957, inst_s15850.g2355, inst_s15850.g2601, inst_s15850.g2602, inst_s15850.g2603, inst_s15850.g2604, inst_s15850.g2605, inst_s15850.g2606, inst_s15850.g2607, inst_s15850.g2608, inst_s15850.g2609, inst_s15850.g2610, inst_s15850.g2611, inst_s15850.g2612, inst_s15850.g2648, inst_s15850.g2986, inst_s15850.g3007, inst_s15850.g3069, inst_s15850.g3327, inst_s15850.g4171, inst_s15850.g4172, inst_s15850.g4173, inst_s15850.g4174, inst_s15850.g4175, inst_s15850.g4176, inst_s15850.g4177, inst_s15850.g4178, inst_s15850.g4179, inst_s15850.g4180, inst_s15850.g4181, inst_s15850.g4191, inst_s15850.g4192, inst_s15850.g4193, inst_s15850.g4194, inst_s15850.g4195, inst_s15850.g4196, inst_s15850.g4197, inst_s15850.g4198, inst_s15850.g4199, inst_s15850.g4200, inst_s15850.g4201, inst_s15850.g4202, inst_s15850.g4203, inst_s15850.g4204, inst_s15850.g4205, inst_s15850.g4206, inst_s15850.g4207, inst_s15850.g4208, inst_s15850.g4209, inst_s15850.g4210, inst_s15850.g4211, inst_s15850.g4212, inst_s15850.g4213, inst_s15850.g4214, inst_s15850.g4215, inst_s15850.g4216, inst_s15850.g4887, inst_s15850.g4888, inst_s15850.g5101, inst_s15850.g5105, inst_s15850.g5658, inst_s15850.g5659, inst_s15850.g5816, inst_s15850.g6253, inst_s15850.g6254, inst_s15850.g6255, inst_s15850.g6256, inst_s15850.g6257, inst_s15850.g6258, inst_s15850.g6259, inst_s15850.g6260, inst_s15850.g6261, inst_s15850.g6262, inst_s15850.g6263, inst_s15850.g6264, inst_s15850.g6265, inst_s15850.g6266, inst_s15850.g6267, inst_s15850.g6268, inst_s15850.g6269, inst_s15850.g6270, inst_s15850.g6271, inst_s15850.g6272, inst_s15850.g6273, inst_s15850.g6274, inst_s15850.g6275, inst_s15850.g6276, inst_s15850.g6277, inst_s15850.g6278, inst_s15850.g6279, inst_s15850.g6280, inst_s15850.g6281, inst_s15850.g6282, inst_s15850.g6283, inst_s15850.g6284, inst_s15850.g6285, inst_s15850.g6842, inst_s15850.g6920, inst_s15850.g6926, inst_s15850.g6932, inst_s15850.g6942, inst_s15850.g6949, inst_s15850.g6955, inst_s15850.g7744, inst_s15850.g8061, inst_s15850.g8062, inst_s15850.g8271, inst_s15850.g8313, inst_s15850.g8316, inst_s15850.g8318, inst_s15850.g8323, inst_s15850.g8328, inst_s15850.g8331, inst_s15850.g8335, inst_s15850.g8340, inst_s15850.g8347, inst_s15850.g8349, inst_s15850.g8352, inst_s15850.g8561, inst_s15850.g8562, inst_s15850.g8563, inst_s15850.g8564, inst_s15850.g8565, inst_s15850.g8566, inst_s15850.g8976, inst_s15850.g8977, inst_s15850.g8978, inst_s15850.g8979, inst_s15850.g8980, inst_s15850.g8981, inst_s15850.g8982, inst_s15850.g8983, inst_s15850.g8984, inst_s15850.g8985, inst_s15850.g8986, inst_s15850.g9451, inst_s15850.g9961, inst_s15850.test_so1, inst_s15850.test_so2, inst_s15850.test_so3, inst_s15850.test_so4, inst_s15850.test_so5, inst_s15850.test_so6, inst_s15850.test_so7, inst_s15850.test_so8, inst_s15850.test_so9, inst_s15850.test_so10, inst_s15850.N599, inst_s15850.g1289, inst_s15850.g1882, inst_s15850.g312, inst_s15850.g452, inst_s15850.g11257, inst_s15850.g123, inst_s15850.g207, inst_s15850.g713, inst_s15850.g1153, inst_s15850.g1744, inst_s15850.g1558, inst_s15850.g695, inst_s15850.g461, inst_s15850.g940, inst_s15850.g976, inst_s15850.g709, inst_s15850.g8432, inst_s15850.g1092, inst_s15850.g1574, inst_s15850.g1864, inst_s15850.g369, inst_s15850.g1580, inst_s15850.g1736, inst_s15850.g1424, inst_s15850.g1737, inst_s15850.g1672, inst_s15850.g1077, inst_s15850.g1231, inst_s15850.g4, inst_s15850.g1104, inst_s15850.g1304, inst_s15850.g7290, inst_s15850.g243, inst_s15850.g1499, inst_s15850.g1444, inst_s15850.g1543, inst_s15850.g315, inst_s15850.g1534, inst_s15850.g622, inst_s15850.g1927, inst_s15850.g1660, inst_s15850.g278, inst_s15850.g1436, inst_s15850.g718, inst_s15850.g8433, inst_s15850.g554, inst_s15850.g496, inst_s15850.g11333, inst_s15850.g981, inst_s15850.g829, inst_s15850.g1095, inst_s15850.g704, inst_s15850.g1265, inst_s15850.g7302, inst_s15850.g1786, inst_s15850.g682, inst_s15850.g8429, inst_s15850.g1296, inst_s15850.g7292, inst_s15850.g327, inst_s15850.g1389, inst_s15850.g1371, inst_s15850.g1956, inst_s15850.g1955, inst_s15850.g1675, inst_s15850.g354, inst_s15850.g113, inst_s15850.g639, inst_s15850.g1684, inst_s15850.g1639, inst_s15850.g1791, inst_s15850.g248, inst_s15850.g1707, inst_s15850.g1759, inst_s15850.g351, inst_s15850.g1604, inst_s15850.g1098, inst_s15850.g932, inst_s15850.g1896, inst_s15850.g8282, inst_s15850.g736, inst_s15850.g8435, inst_s15850.g1019, inst_s15850.g745, inst_s15850.g1419, inst_s15850.g32, inst_s15850.g1086, inst_s15850.g1486, inst_s15850.g1730, inst_s15850.g1504, inst_s15850.g1470, inst_s15850.g822, inst_s15850.g1678, inst_s15850.g174, inst_s15850.g1766, inst_s15850.g1801, inst_s15850.g186, inst_s15850.g959, inst_s15850.g1407, inst_s15850.g1868, inst_s15850.g1718, inst_s15850.g396, inst_s15850.g11265, inst_s15850.g1015, inst_s15850.g1415, inst_s15850.g1227, inst_s15850.g1721, inst_s15850.g284, inst_s15850.g426, inst_s15850.g11256, inst_s15850.g219, inst_s15850.g1360, inst_s15850.g806, inst_s15850.g1428, inst_s15850.g1564, inst_s15850.g1741, inst_s15850.g225, inst_s15850.g281, inst_s15850.g1308, inst_s15850.g611, inst_s15850.g1217, inst_s15850.g1589, inst_s15850.g1466, inst_s15850.g1571, inst_s15850.g1861, inst_s15850.g1448, inst_s15850.g1133, inst_s15850.g1333, inst_s15850.g153, inst_s15850.g962, inst_s15850.g486, inst_s15850.g11331, inst_s15850.g471, inst_s15850.g1397, inst_s15850.g1950, inst_s15850.g8288, inst_s15850.g756, inst_s15850.g755, inst_s15850.g1101, inst_s15850.g549, inst_s15850.g105, inst_s15850.g1669, inst_s15850.g1531, inst_s15850.g1458, inst_s15850.g572, inst_s15850.g1011, inst_s15850.g1411, inst_s15850.g1074, inst_s15850.g444, inst_s15850.g11259, inst_s15850.g1474, inst_s15850.g1080, inst_s15850.g1713, inst_s15850.g333, inst_s15850.g269, inst_s15850.g401, inst_s15850.g11266, inst_s15850.g1857, inst_s15850.g9, inst_s15850.g664, inst_s15850.g965, inst_s15850.g1400, inst_s15850.g309, inst_s15850.g814, inst_s15850.g231, inst_s15850.g557, inst_s15850.g869, inst_s15850.g875, inst_s15850.g1383, inst_s15850.g158, inst_s15850.g627, inst_s15850.g1023, inst_s15850.g259, inst_s15850.g1327, inst_s15850.g654, inst_s15850.g293, inst_s15850.g1346, inst_s15850.g1633, inst_s15850.g1753, inst_s15850.g1508, inst_s15850.g1240, inst_s15850.g7297, inst_s15850.g538, inst_s15850.g11326, inst_s15850.g416, inst_s15850.g11269, inst_s15850.g542, inst_s15850.g11325, inst_s15850.g1681, inst_s15850.g374, inst_s15850.g563, inst_s15850.g1914, inst_s15850.g8284, inst_s15850.g530, inst_s15850.g11328, inst_s15850.g575, inst_s15850.g1936, inst_s15850.g1317, inst_s15850.g1356, inst_s15850.g357, inst_s15850.g386, inst_s15850.g11263, inst_s15850.g1601, inst_s15850.g166, inst_s15850.g501, inst_s15850.g11334, inst_s15850.g262, inst_s15850.g1840, inst_s15850.g318, inst_s15850.g794, inst_s15850.g302, inst_s15850.g342, inst_s15850.g1250, inst_s15850.g7299, inst_s15850.g1163, inst_s15850.g1032, inst_s15850.g1432, inst_s15850.g1453, inst_s15850.g363, inst_s15850.g330, inst_s15850.g1157, inst_s15850.g928, inst_s15850.g261, inst_s15850.g516, inst_s15850.g11337, inst_s15850.g254, inst_s15850.g861, inst_s15850.g1627, inst_s15850.g1292, inst_s15850.g7293, inst_s15850.g290, inst_s15850.g1583, inst_s15850.g466, inst_s15850.g1561, inst_s15850.g1546, inst_s15850.g287, inst_s15850.g560, inst_s15850.g617, inst_s15850.g336, inst_s15850.g456, inst_s15850.g305, inst_s15850.g345, inst_s15850.g8, inst_s15850.g255, inst_s15850.g1945, inst_s15850.g1738, inst_s15850.g1478, inst_s15850.g1690, inst_s15850.g1482, inst_s15850.g1110, inst_s15850.g296, inst_s15850.g1663, inst_s15850.g700, inst_s15850.g8431, inst_s15850.g1762, inst_s15850.g360, inst_s15850.g192, inst_s15850.g1657, inst_s15850.g722, inst_s15850.g566, inst_s15850.g1089, inst_s15850.g1071, inst_s15850.g986, inst_s15850.g971, inst_s15850.g143, inst_s15850.g1814, inst_s15850.g1212, inst_s15850.g1918, inst_s15850.g1822, inst_s15850.g237, inst_s15850.g746, inst_s15850.g1462, inst_s15850.g178, inst_s15850.g366, inst_s15850.g837, inst_s15850.g599, inst_s15850.g1854, inst_s15850.g944, inst_s15850.g1941, inst_s15850.g8287, inst_s15850.g170, inst_s15850.g1520, inst_s15850.g686, inst_s15850.g953, inst_s15850.g1958, inst_s15850.g1765, inst_s15850.g1733, inst_s15850.g7303, inst_s15850.g1610, inst_s15850.g1796, inst_s15850.g1324, inst_s15850.g1540, inst_s15850.g491, inst_s15850.g11332, inst_s15850.g213, inst_s15850.g1781, inst_s15850.g1900, inst_s15850.g1245, inst_s15850.g7298, inst_s15850.g148, inst_s15850.g833, inst_s15850.g1923, inst_s15850.g8285, inst_s15850.g936, inst_s15850.g1314, inst_s15850.g849, inst_s15850.g1336, inst_s15850.g272, inst_s15850.g1806, inst_s15850.g826, inst_s15850.g1887, inst_s15850.g8281, inst_s15850.g968, inst_s15850.g1137, inst_s15850.g1891, inst_s15850.g1255, inst_s15850.g7300, inst_s15850.g257, inst_s15850.g874, inst_s15850.g591, inst_s15850.g731, inst_s15850.g636, inst_s15850.g1218, inst_s15850.g605, inst_s15850.g182, inst_s15850.g950, inst_s15850.g1129, inst_s15850.g857, inst_s15850.g448, inst_s15850.g11258, inst_s15850.g1828, inst_s15850.g1727, inst_s15850.g1592, inst_s15850.g1703, inst_s15850.g1932, inst_s15850.g8286, inst_s15850.g1624, inst_s15850.g440, inst_s15850.g11260, inst_s15850.g476, inst_s15850.g11338, inst_s15850.g119, inst_s15850.g668, inst_s15850.g139, inst_s15850.g1149, inst_s15850.g263, inst_s15850.g818, inst_s15850.g1747, inst_s15850.g802, inst_s15850.g275, inst_s15850.g1524, inst_s15850.g1577, inst_s15850.g810, inst_s15850.g391, inst_s15850.g11264, inst_s15850.g658, inst_s15850.g1386, inst_s15850.g253, inst_s15850.g1125, inst_s15850.g201, inst_s15850.g1280, inst_s15850.g7295, inst_s15850.g1083, inst_s15850.g650, inst_s15850.g1636, inst_s15850.g853, inst_s15850.g421, inst_s15850.g11270, inst_s15850.g956, inst_s15850.g378, inst_s15850.g1756, inst_s15850.g841, inst_s15850.g1027, inst_s15850.g1003, inst_s15850.g1403, inst_s15850.g1145, inst_s15850.g1107, inst_s15850.g1223, inst_s15850.g406, inst_s15850.g11267, inst_s15850.g1811, inst_s15850.g1654, inst_s15850.g197, inst_s15850.g1595, inst_s15850.g1537, inst_s15850.g727, inst_s15850.g8434, inst_s15850.g798, inst_s15850.g481, inst_s15850.g11324, inst_s15850.g1330, inst_s15850.g845, inst_s15850.g1512, inst_s15850.g1490, inst_s15850.g1166, inst_s15850.g348, inst_s15850.g1260, inst_s15850.g7301, inst_s15850.g260, inst_s15850.g131, inst_s15850.g258, inst_s15850.g521, inst_s15850.g11330, inst_s15850.g1318, inst_s15850.g1872, inst_s15850.g677, inst_s15850.g1549, inst_s15850.g947, inst_s15850.g1834, inst_s15850.g1598, inst_s15850.g1121, inst_s15850.g1321, inst_s15850.g506, inst_s15850.g11335, inst_s15850.g546, inst_s15850.g1909, inst_s15850.g1552, inst_s15850.g1687, inst_s15850.g1586, inst_s15850.g324, inst_s15850.g1141, inst_s15850.g1341, inst_s15850.g1710, inst_s15850.g135, inst_s15850.g525, inst_s15850.g11329, inst_s15850.g1607, inst_s15850.g321, inst_s15850.g1275, inst_s15850.g11443, inst_s15850.g1615, inst_s15850.g382, inst_s15850.g266, inst_s15850.g1284, inst_s15850.g7294, inst_s15850.g673, inst_s15850.g8428, inst_s15850.g162, inst_s15850.g411, inst_s15850.g11268, inst_s15850.g431, inst_s15850.g11262, inst_s15850.g1905, inst_s15850.g8283, inst_s15850.g1515, inst_s15850.g1630, inst_s15850.g991, inst_s15850.g1300, inst_s15850.g7291, inst_s15850.g339, inst_s15850.g256, inst_s15850.g1750, inst_s15850.g1440, inst_s15850.g1666, inst_s15850.g1528, inst_s15850.g1351, inst_s15850.g127, inst_s15850.g1618, inst_s15850.g1235, inst_s15850.g7296, inst_s15850.g299, inst_s15850.g435, inst_s15850.g11261, inst_s15850.g1555, inst_s15850.g995, inst_s15850.g1621, inst_s15850.g643, inst_s15850.g1494, inst_s15850.g1567, inst_s15850.g691, inst_s15850.g8430, inst_s15850.g534, inst_s15850.g11327, inst_s15850.g1776, inst_s15850.g569, inst_s15850.g1160, inst_s15850.g1, inst_s15850.g511, inst_s15850.g11336, inst_s15850.g1724, inst_s15850.g12, inst_s15850.g1878, inst_s15850.g4500, inst_s15850.g5529, inst_s15850.g4338, inst_s15850.g8147, inst_s15850.g6551, inst_s15850.g10865, inst_s15850.g8054, inst_s15850.g7709, inst_s15850.g4940, inst_s15850.g6481, inst_s15850.g6529, inst_s15850.g10707, inst_s15850.g6949, inst_s15850.g8940, inst_s15850.g10855, inst_s15850.g6920, inst_s15850.g6907, inst_s15850.g6155, inst_s15850.g6638, inst_s15850.g11647, inst_s15850.g6910, inst_s15850.g6828, inst_s15850.g10800, inst_s15850.g8019, inst_s15850.g6821, inst_s15850.g11478, inst_s15850.g6516, inst_s15850.g8244, inst_s15850.g8631, inst_s15850.g10793, inst_s15850.g5910, inst_s15850.g2478, inst_s15850.g10726, inst_s15850.g6824, inst_s15850.g9961, inst_s15850.g6759, inst_s15850.g6502, inst_s15850.g10797, inst_s15850.g4471, inst_s15850.g10780, inst_s15850.g11625, inst_s15850.g11372, inst_s15850.g10771, inst_s15850.g11293, inst_s15850.g8173, inst_s15850.g6533, inst_s15850.g8245, inst_s15850.g10767, inst_s15850.g6000, inst_s15850.g4490, inst_s15850.g4903, inst_s15850.g10720, inst_s15850.g6934, inst_s15850.g6123, inst_s15850.g6838, inst_s15850.g4905, inst_s15850.g10798, inst_s15850.g10785, inst_s15850.g7204, inst_s15850.g6830, inst_s15850.g8944, inst_s15850.g5543, inst_s15850.g8921, inst_s15850.g6096, inst_s15850.g6942, inst_s15850.g6733, inst_s15850.g6823, inst_s15850.g4890, inst_s15850.g3381, inst_s15850.g10863, inst_s15850.g8039, inst_s15850.g6526, inst_s15850.g10664, inst_s15850.g7189, inst_s15850.g8923, inst_s15850.g5173, inst_s15850.g4264, inst_s15850.g6755, inst_s15850.g11514, inst_s15850.g4506, inst_s15850.g4465, inst_s15850.g6902, inst_s15850.g6015, inst_s15850.g11340, inst_s15850.g6542, inst_s15850.g6507, inst_s15850.g5556, inst_s15850.g8505, inst_s15850.g11641, inst_s15850.g10765, inst_s15850.g11305, inst_s15850.g6126, inst_s15850.g8060, inst_s15850.g7191, inst_s15850.g6469, inst_s15850.g4498, inst_s15850.g6627, inst_s15850.g4893, inst_s15850.g5194, inst_s15850.g6901, inst_s15850.g8043, inst_s15850.g6929, inst_s15850.g8049, inst_s15850.g6786, inst_s15850.g6234, inst_s15850.g10864, inst_s15850.g8984, inst_s15850.g10862, inst_s15850.g10721, inst_s15850.g8051, inst_s15850.g6541, inst_s15850.g10773, inst_s15850.g8193, inst_s15850.g6523, inst_s15850.g5404, inst_s15850.g11393, inst_s15850.g4334, inst_s15850.g6908, inst_s15850.g8768, inst_s15850.g8885, inst_s15850.g6333, inst_s15850.g6045, inst_s15850.g7590, inst_s15850.g6468, inst_s15850.g10782, inst_s15850.g6672, inst_s15850.g6840, inst_s15850.g5914, inst_s15850.g7705, inst_s15850.g6038, inst_s15850.g6471, inst_s15850.g11303, inst_s15850.g10663, inst_s15850.g8920, inst_s15850.g4283, inst_s15850.g4484, inst_s15850.g5396, inst_s15850.g8045, inst_s15850.g7843, inst_s15850.g6932, inst_s15850.g6537, inst_s15850.g4902, inst_s15850.g6080, inst_s15850.g6059, inst_s15850.g4089, inst_s15850.g5126, inst_s15850.g10866, inst_s15850.g11603, inst_s15850.g6332, inst_s15850.g4231, inst_s15850.g11488, inst_s15850.g6955, inst_s15850.g5918, inst_s15850.g6894, inst_s15850.g4076, inst_s15850.g6534, inst_s15850.g6928, inst_s15850.g6926, inst_s15850.g8055, inst_s15850.g11291, inst_s15850.g6833, inst_s15850.g6918, inst_s15850.g6915, inst_s15850.g6911, inst_s15850.g7441, inst_s15850.g5996, inst_s15850.g8047, inst_s15850.g6653, inst_s15850.g6832, inst_s15850.g11481, inst_s15850.g6478, inst_s15850.g6897, inst_s15850.g6042, inst_s15850.g4342, inst_s15850.g4330, inst_s15850.g11609, inst_s15850.g10859, inst_s15850.g6054, inst_s15850.g6508, inst_s15850.g6531, inst_s15850.g8050, inst_s15850.g11376, inst_s15850.g8559, inst_s15850.g7032, inst_s15850.g4293, inst_s15850.g5390, inst_s15850.g8767, inst_s15850.g4480, inst_s15850.g11483, inst_s15850.g5392, inst_s15850.g10776, inst_s15850.g6513, inst_s15850.g9272, inst_s15850.g10898, inst_s15850.g8052, inst_s15850.g4325, inst_s15850.g8766, inst_s15850.g6205, inst_s15850.g8820, inst_s15850.g9124, inst_s15850.g6839, inst_s15850.g6522, inst_s15850.g10936, inst_s15850.g11320, inst_s15850.g6841, inst_s15850.g8769, inst_s15850.g6224, inst_s15850.g11349, inst_s15850.g6470, inst_s15850.g5755, inst_s15850.g6515, inst_s15850.g10791, inst_s15850.g7632, inst_s15850.g11485, inst_s15850.g6331, inst_s15850.g8053, inst_s15850.g5763, inst_s15850.g6480, inst_s15850.g6795, inst_s15850.g8194, inst_s15850.g8938, inst_s15850.g4238, inst_s15850.g8775, inst_s15850.g4891, inst_s15850.g11290, inst_s15850.g6501, inst_s15850.g6334, inst_s15850.g10719, inst_s15850.g4274, inst_s15850.g8765, inst_s15850.g6916, inst_s15850.g11308, inst_s15850.g10784, inst_s15850.g6820, inst_s15850.g4340, inst_s15850.g6922, inst_s15850.g6747, inst_s15850.g11391, inst_s15850.g8649, inst_s15850.g9555, inst_s15850.g6071, inst_s15850.g10858, inst_s15850.g8926, inst_s15850.g4239, inst_s15850.g11602, inst_s15850.g8041, inst_s15850.g8922, inst_s15850.g5536, inst_s15850.g11605, inst_s15850.g8048, inst_s15850.g6528, inst_s15850.g6524, inst_s15850.g7219, inst_s15850.g8046, inst_s15850.g11482, inst_s15850.g4477, inst_s15850.g6923, inst_s15850.g4255, inst_s15850.g8937, inst_s15850.g6538, inst_s15850.g11306, inst_s15850.g7183, inst_s15850.g6895, inst_s15850.g6179, inst_s15850.g9721, inst_s15850.g8776, inst_s15850.g6827, inst_s15850.g4309, inst_s15850.g7244, inst_s15850.g7586, inst_s15850.g7930, inst_s15850.g11300, inst_s15850.g10718, inst_s15850.g5445, inst_s15850.g6088, inst_s15850.g6679, inst_s15850.g11636, inst_s15850.g9266, inst_s15850.g11608, inst_s15850.g8059, inst_s15850.g8771, inst_s15850.g6035, inst_s15850.g6198, inst_s15850.g8973, inst_s15850.g6834, inst_s15850.g5148, inst_s15850.g7134, inst_s15850.g10795, inst_s15850.g10770, inst_s15850.g8773, inst_s15850.g3462, inst_s15850.g7143, inst_s15850.g8939, inst_s15850.g8772, inst_s15850.g6093, inst_s15850.g6500, inst_s15850.g8777, inst_s15850.g6244, inst_s15850.g11640, inst_s15850.g11487, inst_s15850.g9110, inst_s15850.g11380, inst_s15850.g9269, inst_s15850.g11314, inst_s15850.g9150, inst_s15850.g11298, inst_s15850.g7202, inst_s15850.g6819, inst_s15850.g6243, inst_s15850.g6514, inst_s15850.g6983, inst_s15850.g4473, inst_s15850.g8040, inst_s15850.g6900, inst_s15850.g8042, inst_s15850.g6546, inst_s15850.g5770, inst_s15850.g8889, inst_s15850.g10711, inst_s15850.g11312, inst_s15850.g6479, inst_s15850.g5849, inst_s15850.g6656, inst_s15850.g6906, inst_s15850.g10717, inst_s15850.g8770, inst_s15850.g6392, inst_s15850.g6621, inst_s15850.g11610, inst_s15850.g11604, inst_s15850.g11486, inst_s15850.g7581, inst_s15850.g10799, inst_s15850.g6439, inst_s15850.g7133, inst_s15850.g8044, inst_s15850.g8254, inst_s15850.g11607, inst_s15850.g6193, inst_s15850.g4904, inst_s15850.g11292, inst_s15850.g6822, inst_s15850.g6912, inst_s15850.g6898, inst_s15850.g5421, inst_s15850.g6924, inst_s15850.g11310, inst_s15850.g11294, inst_s15850.g6026, inst_s15850.g8024, inst_s15850.g8945, inst_s15850.g6525, inst_s15850.g5083, inst_s15850.g7541, inst_s15850.g10860, inst_s15850.g11579, inst_s15850.g11639, inst_s15850.g6826, inst_s15850.g7626, inst_s15850.g6829, inst_s15850.g7660, inst_s15850.g10722, inst_s15850.g8887, inst_s15850.g11484, inst_s15850.g6002, inst_s15850.g11606, inst_s15850.g6757, inst_s15850.g6216, inst_s15850.g8941, inst_s15850.g4892, inst_s15850.g6930, inst_s15850.g8250, inst_s15850.g6049, inst_s15850.g8943, inst_s15850.g10861, inst_s15850.g8779, inst_s15850.g6180, inst_s15850.g8774, inst_s15850.g8260, inst_s15850.g6099, inst_s15850.g6831, inst_s15850.g6068, inst_s15850.g7137, inst_s15850.g6545, inst_s15850.g7257, inst_s15850.g6909, inst_s15850.g8384, inst_s15850.g11392, inst_s15850.g6506, inst_s15850.g8883, inst_s15850.g6728, inst_s15850.g10724, inst_s15850.g4556, inst_s15850.DFF_121_n1, inst_s15850.DFF_122_n1, inst_s15850.DFF_126_n1, inst_s15850.DFF_136_n1, inst_s15850.DFF_157_n1, inst_s15850.DFF_168_n1, inst_s15850.DFF_194_n1, inst_s15850.DFF_228_n1, inst_s15850.g8271, inst_s15850.DFF_242_n1, inst_s15850.DFF_275_n1, inst_s15850.DFF_311_n1, inst_s15850.DFF_319_n1, inst_s15850.DFF_330_n1, inst_s15850.DFF_336_n1, inst_s15850.DFF_350_n1, inst_s15850.DFF_384_n1, inst_s15850.DFF_385_n1, inst_s15850.DFF_436_n1, inst_s15850.DFF_441_n1, inst_s15850.DFF_445_n1, inst_s15850.DFF_452_n1, inst_s15850.DFF_489_n1, inst_s15850.n517, inst_s15850.n518, inst_s15850.n519, inst_s15850.n520, inst_s15850.n521, inst_s15850.n522, inst_s15850.n524, inst_s15850.n526, inst_s15850.n527, inst_s15850.n528, inst_s15850.n529, inst_s15850.n530, inst_s15850.n532, inst_s15850.n533, inst_s15850.n534, inst_s15850.n535, inst_s15850.n536, inst_s15850.n537, inst_s15850.n538, inst_s15850.n539, inst_s15850.n540, inst_s15850.n542, inst_s15850.n544, inst_s15850.n545, inst_s15850.n546, inst_s15850.n547, inst_s15850.n548, inst_s15850.n549, inst_s15850.n550, inst_s15850.n551, inst_s15850.n552, inst_s15850.n553, inst_s15850.n554, inst_s15850.n555, inst_s15850.n556, inst_s15850.n557, inst_s15850.n560, inst_s15850.n561, inst_s15850.n562, inst_s15850.n563, inst_s15850.n564, inst_s15850.n565, inst_s15850.n566, inst_s15850.n567, inst_s15850.n568, inst_s15850.n569, inst_s15850.n572, inst_s15850.n573, inst_s15850.n574, inst_s15850.n575, inst_s15850.n576, inst_s15850.n577, inst_s15850.n578, inst_s15850.n579, inst_s15850.n580, inst_s15850.n581, inst_s15850.n583, inst_s15850.n592, inst_s15850.n594, inst_s15850.n595, inst_s15850.n596, inst_s15850.n597, inst_s15850.n598, inst_s15850.n599, inst_s15850.n600, inst_s15850.n602, inst_s15850.n603, inst_s15850.n604, inst_s15850.n605, inst_s15850.n606, inst_s15850.n607, inst_s15850.n609, inst_s15850.n610, inst_s15850.n611, inst_s15850.n612, inst_s15850.n614, inst_s15850.n616, inst_s15850.n617, inst_s15850.n619, inst_s15850.n620, inst_s15850.n621, inst_s15850.n622, inst_s15850.n623, inst_s15850.n624, inst_s15850.n625, inst_s15850.n627, inst_s15850.n629, inst_s15850.n630, inst_s15850.n631, inst_s15850.n632, inst_s15850.n633, inst_s15850.n634, inst_s15850.n643, inst_s15850.n644, inst_s15850.n645, inst_s15850.n646, inst_s15850.n647, inst_s15850.n648, inst_s15850.n649, inst_s15850.n650, inst_s15850.n651, inst_s15850.n661, inst_s15850.n662, inst_s15850.n665, inst_s15850.n667, inst_s15850.n668, inst_s15850.n674, inst_s15850.n675, inst_s15850.n685, inst_s15850.n687, inst_s15850.n711, inst_s15850.n712, inst_s15850.n713, inst_s15850.n715, inst_s15850.n717, inst_s15850.n718, inst_s15850.n719, inst_s15850.n720, inst_s15850.n721, inst_s15850.n725, inst_s15850.n744, inst_s15850.n793, inst_s15850.n794, inst_s15850.n795, inst_s15850.n796, inst_s15850.n797, inst_s15850.n798, inst_s15850.n799, inst_s15850.n800, inst_s15850.n801, inst_s15850.n802, inst_s15850.n803, inst_s15850.n804, inst_s15850.n805, inst_s15850.n806, inst_s15850.n807, inst_s15850.n808, inst_s15850.n809, inst_s15850.n810, inst_s15850.n811, inst_s15850.n812, inst_s15850.n813, inst_s15850.n814, inst_s15850.n815, inst_s15850.n816, inst_s15850.n817, inst_s15850.n818, inst_s15850.n819, inst_s15850.n820, inst_s15850.n821, inst_s15850.n822, inst_s15850.n823, inst_s15850.n824, inst_s15850.n825, inst_s15850.n826, inst_s15850.n827, inst_s15850.n828, inst_s15850.n829, inst_s15850.n830, inst_s15850.n831, inst_s15850.n832, inst_s15850.n833, inst_s15850.n834, inst_s15850.n835, inst_s15850.n836, inst_s15850.n837, inst_s15850.n838, inst_s15850.n839, inst_s15850.n840, inst_s15850.n841, inst_s15850.n842, inst_s15850.n843, inst_s15850.n844, inst_s15850.n845, inst_s15850.n846, inst_s15850.n847, inst_s15850.n848, inst_s15850.n849, inst_s15850.n850, inst_s15850.n851, inst_s15850.n852, inst_s15850.n853, inst_s15850.n854, inst_s15850.n855, inst_s15850.n856, inst_s15850.n857, inst_s15850.n858, inst_s15850.n859, inst_s15850.n860, inst_s15850.n861, inst_s15850.n862, inst_s15850.n863, inst_s15850.n864, inst_s15850.n865, inst_s15850.n866, inst_s15850.n867, inst_s15850.n868, inst_s15850.n869, inst_s15850.n870, inst_s15850.n871, inst_s15850.n872, inst_s15850.n873, inst_s15850.n874, inst_s15850.n875, inst_s15850.n876, inst_s15850.n877, inst_s15850.n878, inst_s15850.n879, inst_s15850.n880, inst_s15850.n881, inst_s15850.n882, inst_s15850.n883, inst_s15850.n884, inst_s15850.n885, inst_s15850.n886, inst_s15850.n887, inst_s15850.n888, inst_s15850.n889, inst_s15850.n890, inst_s15850.n891, inst_s15850.n892, inst_s15850.n893, inst_s15850.n894, inst_s15850.n895, inst_s15850.n896, inst_s15850.n897, inst_s15850.n898, inst_s15850.n899, inst_s15850.n900, inst_s15850.n901, inst_s15850.n902, inst_s15850.n903, inst_s15850.n904, inst_s15850.n905, inst_s15850.n906, inst_s15850.n907, inst_s15850.n908, inst_s15850.n909, inst_s15850.n910, inst_s15850.n911, inst_s15850.n912, inst_s15850.n913, inst_s15850.n914, inst_s15850.n915, inst_s15850.n916, inst_s15850.n917, inst_s15850.n918, inst_s15850.n919, inst_s15850.n920, inst_s15850.n921, inst_s15850.n922, inst_s15850.n923, inst_s15850.n924, inst_s15850.n925, inst_s15850.n926, inst_s15850.n927, inst_s15850.n928, inst_s15850.n929, inst_s15850.n930, inst_s15850.n931, inst_s15850.n932, inst_s15850.n933, inst_s15850.n934, inst_s15850.n935, inst_s15850.n936, inst_s15850.n937, inst_s15850.n938, inst_s15850.n939, inst_s15850.n940, inst_s15850.n941, inst_s15850.n942, inst_s15850.n943, inst_s15850.n944, inst_s15850.n945, inst_s15850.n946, inst_s15850.n947, inst_s15850.n948, inst_s15850.n949, inst_s15850.n950, inst_s15850.n951, inst_s15850.n952, inst_s15850.n953, inst_s15850.n954, inst_s15850.n955, inst_s15850.n956, inst_s15850.n957, inst_s15850.n958, inst_s15850.n959, inst_s15850.n960, inst_s15850.n961, inst_s15850.n962, inst_s15850.n963, inst_s15850.n964, inst_s15850.n965, inst_s15850.n966, inst_s15850.n967, inst_s15850.n968, inst_s15850.n969, inst_s15850.n970, inst_s15850.n971, inst_s15850.n972, inst_s15850.n973, inst_s15850.n974, inst_s15850.n975, inst_s15850.n976, inst_s15850.n977, inst_s15850.n978, inst_s15850.n979, inst_s15850.n980, inst_s15850.n981, inst_s15850.n982, inst_s15850.n983, inst_s15850.n984, inst_s15850.n985, inst_s15850.n986, inst_s15850.n987, inst_s15850.n988, inst_s15850.n989, inst_s15850.n990, inst_s15850.n991, inst_s15850.n992, inst_s15850.n993, inst_s15850.n994, inst_s15850.n995, inst_s15850.n996, inst_s15850.n997, inst_s15850.n998, inst_s15850.n999, inst_s15850.n1000, inst_s15850.n1001, inst_s15850.n1002, inst_s15850.n1003, inst_s15850.n1004, inst_s15850.n1005, inst_s15850.n1006, inst_s15850.n1007, inst_s15850.n1008, inst_s15850.n1009, inst_s15850.n1010, inst_s15850.n1011, inst_s15850.n1012, inst_s15850.n1013, inst_s15850.n1014, inst_s15850.n1015, inst_s15850.n1016, inst_s15850.n1017, inst_s15850.n1018, inst_s15850.n1019, inst_s15850.n1020, inst_s15850.n1021, inst_s15850.n1022, inst_s15850.n1023, inst_s15850.n1024, inst_s15850.n1025, inst_s15850.n1026, inst_s15850.n1027, inst_s15850.n1028, inst_s15850.n1029, inst_s15850.n1030, inst_s15850.n1031, inst_s15850.n1032, inst_s15850.n1033, inst_s15850.n1034, inst_s15850.n1035, inst_s15850.n1036, inst_s15850.n1037, inst_s15850.n1038, inst_s15850.n1039, inst_s15850.n1040, inst_s15850.n1041, inst_s15850.n1042, inst_s15850.n1043, inst_s15850.n1044, inst_s15850.n1045, inst_s15850.n1046, inst_s15850.n1047, inst_s15850.n1048, inst_s15850.n1049, inst_s15850.n1050, inst_s15850.n1051, inst_s15850.n1052, inst_s15850.n1053, inst_s15850.n1054, inst_s15850.n1055, inst_s15850.n1056, inst_s15850.n1057, inst_s15850.n1058, inst_s15850.n1059, inst_s15850.n1060, inst_s15850.n1061, inst_s15850.n1062, inst_s15850.n1063, inst_s15850.n1064, inst_s15850.n1065, inst_s15850.n1066, inst_s15850.n1067, inst_s15850.n1068, inst_s15850.n1069, inst_s15850.n1070, inst_s15850.n1071, inst_s15850.n1072, inst_s15850.n1073, inst_s15850.n1074, inst_s15850.n1075, inst_s15850.n1076, inst_s15850.n1077, inst_s15850.n1078, inst_s15850.n1079, inst_s15850.n1080, inst_s15850.n1081, inst_s15850.n1082, inst_s15850.n1083, inst_s15850.n1084, inst_s15850.n1085, inst_s15850.n1086, inst_s15850.n1087, inst_s15850.n1088, inst_s15850.n1089, inst_s15850.n1090, inst_s15850.n1091, inst_s15850.n1092, inst_s15850.n1093, inst_s15850.n1094, inst_s15850.n1095, inst_s15850.n1096, inst_s15850.n1097, inst_s15850.n1098, inst_s15850.n1099, inst_s15850.n1100, inst_s15850.n1101, inst_s15850.n1102, inst_s15850.n1103, inst_s15850.n1104, inst_s15850.n1105, inst_s15850.n1106, inst_s15850.n1107, inst_s15850.n1108, inst_s15850.n1109, inst_s15850.n1110, inst_s15850.n1111, inst_s15850.n1112, inst_s15850.n1113, inst_s15850.n1114, inst_s15850.n1115, inst_s15850.n1116, inst_s15850.n1117, inst_s15850.n1118, inst_s15850.n1119, inst_s15850.n1120, inst_s15850.n1122, inst_s15850.n1123, inst_s15850.n1124, inst_s15850.n1125, inst_s15850.n1126, inst_s15850.n1127, inst_s15850.n1128, inst_s15850.n1129, inst_s15850.n1130, inst_s15850.n1131, inst_s15850.n1132, inst_s15850.n1133, inst_s15850.n1134, inst_s15850.n1135, inst_s15850.n1136, inst_s15850.n1137, inst_s15850.n1138, inst_s15850.n1139, inst_s15850.n1140, inst_s15850.n1141, inst_s15850.n1142, inst_s15850.n1143, inst_s15850.n1144, inst_s15850.n1145, inst_s15850.n1146, inst_s15850.n1147, inst_s15850.n1148, inst_s15850.n1149, inst_s15850.n1150, inst_s15850.n1151, inst_s15850.n1152, inst_s15850.n1153, inst_s15850.n1154, inst_s15850.n1155, inst_s15850.n1156, inst_s15850.n1157, inst_s15850.n1158, inst_s15850.n1159, inst_s15850.n1160, inst_s15850.n1161, inst_s15850.n1162, inst_s15850.n1163, inst_s15850.n1164, inst_s15850.n1165, inst_s15850.n1166, inst_s15850.n1167, inst_s15850.n1168, inst_s15850.n1169, inst_s15850.n1170, inst_s15850.n1171, inst_s15850.n1172, inst_s15850.n1173, inst_s15850.n1174, inst_s15850.n1175, inst_s15850.n1176, inst_s15850.n1177, inst_s15850.n1178, inst_s15850.n1179, inst_s15850.n1180, inst_s15850.n1181, inst_s15850.n1182, inst_s15850.n1183, inst_s15850.n1184, inst_s15850.n1185, inst_s15850.n1186, inst_s15850.n1187, inst_s15850.n1188, inst_s15850.n1189, inst_s15850.n1190, inst_s15850.n1191, inst_s15850.n1192, inst_s15850.n1193, inst_s15850.n1195, inst_s15850.n1196, inst_s15850.n1197, inst_s15850.n1198, inst_s15850.n1199, inst_s15850.n1200, inst_s15850.n1201, inst_s15850.n1202, inst_s15850.n1203, inst_s15850.n1204, inst_s15850.n1205, inst_s15850.n1206, inst_s15850.n1207, inst_s15850.n1208, inst_s15850.n1209, inst_s15850.n1210, inst_s15850.n1211, inst_s15850.n1212, inst_s15850.n1213, inst_s15850.n1214, inst_s15850.n1215, inst_s15850.n1216, inst_s15850.n1217, inst_s15850.n1218, inst_s15850.n1219, inst_s15850.n1220, inst_s15850.n1221, inst_s15850.n1222, inst_s15850.n1223, inst_s15850.n1224, inst_s15850.n1225, inst_s15850.n1226, inst_s15850.n1227, inst_s15850.n1228, inst_s15850.n1229, inst_s15850.n1230, inst_s15850.n1231, inst_s15850.n1232, inst_s15850.n1233, inst_s15850.n1234, inst_s15850.n1235, inst_s15850.n1236, inst_s15850.n1237, inst_s15850.n1238, inst_s15850.n1239, inst_s15850.n1240, inst_s15850.n1241, inst_s15850.n1243, inst_s15850.n1244, inst_s15850.n1245, inst_s15850.n1246, inst_s15850.n1247, inst_s15850.n1248, inst_s15850.n1249, inst_s15850.n1250, inst_s15850.n1251, inst_s15850.n1252, inst_s15850.n1253, inst_s15850.n1254, inst_s15850.n1255, inst_s15850.n1256, inst_s15850.n1257, inst_s15850.n1258, inst_s15850.n1259, inst_s15850.n1260, inst_s15850.n1261, inst_s15850.n1262, inst_s15850.n1263, inst_s15850.n1264, inst_s15850.n1265, inst_s15850.n1266, inst_s15850.n1267, inst_s15850.n1268, inst_s15850.n1269, inst_s15850.n1270, inst_s15850.n1271, inst_s15850.n1272, inst_s15850.n1273, inst_s15850.n1274, inst_s15850.n1275, inst_s15850.n1276, inst_s15850.n1277, inst_s15850.n1278, inst_s15850.n1279, inst_s15850.n1280, inst_s15850.n1281, inst_s15850.n1282, inst_s15850.n1283, inst_s15850.n1284, inst_s15850.n1285, inst_s15850.n1286, inst_s15850.n1287, inst_s15850.n1288, inst_s15850.n1289, inst_s15850.n1290, inst_s15850.n1291, inst_s15850.n1292, inst_s15850.n1293, inst_s15850.n1294, inst_s15850.n1295, inst_s15850.n1296, inst_s15850.n1297, inst_s15850.n1298, inst_s15850.n1299, inst_s15850.n1300, inst_s15850.n1301, inst_s15850.n1302, inst_s15850.n1303, inst_s15850.n1304, inst_s15850.n1305, inst_s15850.n1306, inst_s15850.n1307, inst_s15850.n1308, inst_s15850.n1309, inst_s15850.n1310, inst_s15850.n1311, inst_s15850.n1312, inst_s15850.n1313, inst_s15850.n1314, inst_s15850.n1315, inst_s15850.n1316, inst_s15850.n1317, inst_s15850.n1318, inst_s15850.n1319, inst_s15850.n1320, inst_s15850.n1321, inst_s15850.n1322, inst_s15850.n1323, inst_s15850.n1324, inst_s15850.n1325, inst_s15850.n1326, inst_s15850.n1328, inst_s15850.n1329, inst_s15850.n1330, inst_s15850.n1331, inst_s15850.n1332, inst_s15850.n1333, inst_s15850.n1334, inst_s15850.n1335, inst_s15850.n1336, inst_s15850.n1337, inst_s15850.n1338, inst_s15850.n1339, inst_s15850.n1340, inst_s15850.n1341, inst_s15850.n1342, inst_s15850.n1343, inst_s15850.n1344, inst_s15850.n1345, inst_s15850.n1346, inst_s15850.n1347, inst_s15850.n1348, inst_s15850.n1349, inst_s15850.n1350, inst_s15850.n1351, inst_s15850.n1352, inst_s15850.n1353, inst_s15850.n1354, inst_s15850.n1355, inst_s15850.n1356, inst_s15850.n1357, inst_s15850.n1358, inst_s15850.n1359, inst_s15850.n1360, inst_s15850.n1361, inst_s15850.n1362, inst_s15850.n1363, inst_s15850.n1364, inst_s15850.n1365, inst_s15850.n1366, inst_s15850.n1367, inst_s15850.n1368, inst_s15850.n1369, inst_s15850.n1370, inst_s15850.n1371, inst_s15850.n1372, inst_s15850.n1373, inst_s15850.n1374, inst_s15850.n1375, inst_s15850.n1376, inst_s15850.n1377, inst_s15850.n1378, inst_s15850.n1379, inst_s15850.n1380, inst_s15850.n1381, inst_s15850.n1382, inst_s15850.n1383, inst_s15850.n1384, inst_s15850.n1385, inst_s15850.n1386, inst_s15850.n1387, inst_s15850.n1388, inst_s15850.n1389, inst_s15850.n1390, inst_s15850.n1391, inst_s15850.n1392, inst_s15850.n1393, inst_s15850.n1394, inst_s15850.n1395, inst_s15850.n1396, inst_s15850.n1397, inst_s15850.n1398, inst_s15850.n1399, inst_s15850.n1402, inst_s15850.n1403, inst_s15850.n1404, inst_s15850.n1405, inst_s15850.n1406, inst_s15850.n1407, inst_s15850.n1408, inst_s15850.n1409, inst_s15850.n1410, inst_s15850.n1411, inst_s15850.n1412, inst_s15850.n1413, inst_s15850.n1414, inst_s15850.n1415, inst_s15850.n1416, inst_s15850.n1417, inst_s15850.n1418, inst_s15850.n1419, inst_s15850.n1420, inst_s15850.n1421, inst_s15850.n1422, inst_s15850.n1423, inst_s15850.n1424, inst_s15850.n1425, inst_s15850.n1426, inst_s15850.n1427, inst_s15850.n1428, inst_s15850.n1429, inst_s15850.n1430, inst_s15850.n1431, inst_s15850.n1432, inst_s15850.n1433, inst_s15850.n1434, inst_s15850.n1436, inst_s15850.n1437, inst_s15850.n1438, inst_s15850.n1439, inst_s15850.n1440, inst_s15850.n1441, inst_s15850.n1442, inst_s15850.n1443, inst_s15850.n1444, inst_s15850.n1445, inst_s15850.n1446, inst_s15850.n1447, inst_s15850.n1448, inst_s15850.n1449, inst_s15850.n1450, inst_s15850.n1451, inst_s15850.n1452, inst_s15850.n1453, inst_s15850.n1454, inst_s15850.n1455, inst_s15850.n1459, inst_s15850.n1461, inst_s15850.n1462, inst_s15850.n1463, inst_s15850.n1464, inst_s15850.n1465, inst_s15850.n1466, inst_s15850.n1467, inst_s15850.n1468, inst_s15850.n1469, inst_s15850.n1470, inst_s15850.n1471, inst_s15850.n1472, inst_s15850.n1473, inst_s15850.n1474, inst_s15850.n1475, inst_s15850.n1476, inst_s15850.n1477, inst_s15850.n1478, inst_s15850.n1479, inst_s15850.n1480, inst_s15850.n1481, inst_s15850.n1482, inst_s15850.n1483, inst_s15850.n1484, inst_s15850.n1485, inst_s15850.n1486, inst_s15850.n1487, inst_s15850.n1488, inst_s15850.n1489, inst_s15850.n1490, inst_s15850.n1491, inst_s15850.n1492, inst_s15850.n1493, inst_s15850.n1494, inst_s15850.n1495, inst_s15850.n1496, inst_s15850.n1497, inst_s15850.n1498, inst_s15850.n1499, inst_s15850.n1500, inst_s15850.n1501, inst_s15850.n1502, inst_s15850.n1503, inst_s15850.n1504, inst_s15850.n1505, inst_s15850.n1506, inst_s15850.n1507, inst_s15850.n1508, inst_s15850.n1509, inst_s15850.n1510, inst_s15850.n1511, inst_s15850.n1512, inst_s15850.n1513, inst_s15850.n1514, inst_s15850.n1515, inst_s15850.n1516, inst_s15850.n1517, inst_s15850.n1518, inst_s15850.n1519, inst_s15850.n1520, inst_s15850.n1521, inst_s15850.n1522, inst_s15850.n1523, inst_s15850.n1524, inst_s15850.n1525, inst_s15850.n1526, inst_s15850.n1527, inst_s15850.n1528, inst_s15850.n1529, inst_s15850.n1530, inst_s15850.n1531, inst_s15850.n1532, inst_s15850.n1533, inst_s15850.n1534, inst_s15850.n1535, inst_s15850.n1536, inst_s15850.n1537, inst_s15850.n1538, inst_s15850.n1539, inst_s15850.n1540, inst_s15850.n1541, inst_s15850.n1542, inst_s15850.n1543, inst_s15850.n1544, inst_s15850.n1545, inst_s15850.n1546, inst_s15850.n1547, inst_s15850.n1548, inst_s15850.n1549, inst_s15850.n1550, inst_s15850.n1551, inst_s15850.n1552, inst_s15850.n1553, inst_s15850.n1554, inst_s15850.n1555, inst_s15850.n1556, inst_s15850.n1557, inst_s15850.n1558, inst_s15850.n1559, inst_s15850.n1560, inst_s15850.n1561, inst_s15850.n1562, inst_s15850.n1563, inst_s15850.n1564, inst_s15850.n1565, inst_s15850.n1566, inst_s15850.n1567, inst_s15850.n1568, inst_s15850.n1569, inst_s15850.n1570, inst_s15850.n1571, inst_s15850.n1572, inst_s15850.n1573, inst_s15850.n1574, inst_s15850.n1575, inst_s15850.n1576, inst_s15850.n1577, inst_s15850.n1578, inst_s15850.n1579, inst_s15850.n1580, inst_s15850.n1581, inst_s15850.n1583, inst_s15850.n1585, inst_s15850.n1586, inst_s15850.n1587, inst_s15850.n1588, inst_s15850.n1590, inst_s15850.n1591, inst_s15850.n1592, inst_s15850.n1593, inst_s15850.n1594, inst_s15850.n1595, inst_s15850.n1596, inst_s15850.n1597, inst_s15850.n1598, inst_s15850.n1599, inst_s15850.n1600, inst_s15850.n1601, inst_s15850.n1602, inst_s15850.n1603, inst_s15850.n1604, inst_s15850.n1605, inst_s15850.n1606, inst_s15850.n1607, inst_s15850.n1608, inst_s15850.n1609, inst_s15850.n1610, inst_s15850.n1611, inst_s15850.n1612, inst_s15850.n1613, inst_s15850.n1614, inst_s15850.n1615, inst_s15850.n1616, inst_s15850.n1617, inst_s15850.n1618, inst_s15850.n1619, inst_s15850.n1620, inst_s15850.n1621, inst_s15850.n1622, inst_s15850.n1623, inst_s15850.n1624, inst_s15850.n1625, inst_s15850.n1626, inst_s15850.n1627, inst_s15850.n1628, inst_s15850.n1629, inst_s15850.n1630, inst_s15850.n1631, inst_s15850.n1632, inst_s15850.n1633, inst_s15850.n1634, inst_s15850.n1635, inst_s15850.n1636, inst_s15850.n1637, inst_s15850.n1638, inst_s15850.n1639, inst_s15850.n1640, inst_s15850.n1641, inst_s15850.n1642, inst_s15850.n1643, inst_s15850.n1644, inst_s15850.n1645, inst_s15850.n1646, inst_s15850.n1647, inst_s15850.n1648, inst_s15850.n1649, inst_s15850.n1650, inst_s15850.n1651, inst_s15850.n1652, inst_s15850.n1653, inst_s15850.n1654, inst_s15850.n1655, inst_s15850.n1656, inst_s15850.n1657, inst_s15850.n1658, inst_s15850.n1659, inst_s15850.n1660, inst_s15850.n1661, inst_s15850.n1662, inst_s15850.n1663, inst_s15850.n1664, inst_s15850.n1665, inst_s15850.n1666, inst_s15850.n1667, inst_s15850.n1668, inst_s15850.n1669, inst_s15850.n1670, inst_s15850.n1671, inst_s15850.n1672, inst_s15850.n1673, inst_s15850.n1674, inst_s15850.n1675, inst_s15850.n1676, inst_s15850.n1677, inst_s15850.n1678, inst_s15850.n1679, inst_s15850.n1680, inst_s15850.n1681, inst_s15850.n1682, inst_s15850.n1683, inst_s15850.n1684, inst_s15850.n1685, inst_s15850.n1686, inst_s15850.n1687, inst_s15850.n1688, inst_s15850.n1689, inst_s15850.n1690, inst_s15850.n1691, inst_s15850.n1692, inst_s15850.n1693, inst_s15850.n1694, inst_s15850.n1695, inst_s15850.n1696, inst_s15850.n1697, inst_s15850.n1698, inst_s15850.n1699, inst_s15850.n1700, inst_s15850.n1701, inst_s15850.n1702, inst_s15850.n1703, inst_s15850.n1704, inst_s15850.n1705, inst_s15850.n1706, inst_s15850.n1707, inst_s15850.n1708, inst_s15850.n1709, inst_s15850.n1710, inst_s15850.n1711, inst_s15850.n1712, inst_s15850.n1713, inst_s15850.n1714, inst_s15850.n1715, inst_s15850.n1716, inst_s15850.n1717, inst_s15850.n1718, inst_s15850.n1719, inst_s15850.n1720, inst_s15850.n1721, inst_s15850.n1722, inst_s15850.n1723, inst_s15850.n1724, inst_s15850.n1725, inst_s15850.n1727, inst_s15850.n1729, inst_s15850.n1731, inst_s15850.n1733, inst_s15850.n1735, inst_s15850.n1737, inst_s15850.n1739, inst_s15850.n1741, inst_s15850.n1743, inst_s15850.n1745, inst_s15850.n1747, inst_s15850.n1749, inst_s15850.n1751, inst_s15850.n1753, inst_s15850.n1755, inst_s15850.n1757, inst_s15850.n1759, inst_s15850.n1761, inst_s15850.n1763, inst_s15850.n1765, inst_s15850.n1767, inst_s15850.n1769, inst_s15850.n1771, inst_s15850.n1773, inst_s15850.n1775, inst_s15850.n1777, inst_s15850.n1779, inst_s15850.n1781, inst_s15850.n1783, inst_s15850.n1785, inst_s15850.n1787, inst_s15850.n1789, inst_s15850.n1791, inst_s15850.n1793, inst_s15850.n1795, inst_s15850.n1797, inst_s15850.n1799, inst_s15850.n1801, inst_s15850.n1803, inst_s15850.n1805, inst_s15850.n1807, inst_s15850.n1809, inst_s15850.n1811, inst_s15850.n1813, inst_s15850.n1815, inst_s15850.n1817, inst_s15850.n1819, inst_s15850.n1821, inst_s15850.n1823, inst_s15850.n1825, inst_s15850.n1827, inst_s15850.n1829, inst_s15850.n1831, inst_s15850.n1833, inst_s15850.n1835, inst_s15850.n1837, inst_s15850.g5105, inst_s15850.n1839, inst_s15850.g5101, inst_s15850.n1841, inst_s15850.n1843, inst_s15850.n1845, inst_s15850.n1847, inst_s15850.n1849, inst_s15850.n1851, inst_s15850.n1853, inst_s15850.n1854, inst_s15850.n1855, inst_s15850.n1856, inst_s15850.n1857, inst_s15850.n1858, inst_s15850.n1859, inst_s15850.n1860, inst_s15850.n1861, inst_s15850.n1862, inst_s15850.n1863, inst_s15850.n1864, inst_s15850.n1865, inst_s15850.n1866, inst_s15850.n1867, inst_s15850.n1868, inst_s15850.n1869, inst_s15850.n1870, inst_s15850.n1871, inst_s15850.n1872, inst_s15850.n1873, inst_s15850.n1874, inst_s15850.n1875, inst_s15850.n1876, inst_s15850.n1877, inst_s15850.n1878, inst_s15850.n1880, inst_s15850.n1881, inst_s15850.n1882, inst_s15850.n1883, inst_s15850.n1884, inst_s15850.n1885, inst_s15850.n1886, inst_s15850.n1887, inst_s15850.n1888, inst_s15850.n1889, inst_s15850.n1890, inst_s15850.n1891, inst_s15850.n1892, inst_s15850.n1893, inst_s15850.n1894, inst_s15850.n1895, inst_s15850.n1896, inst_s15850.n1897, inst_s15850.n1898, inst_s15850.n1899, inst_s15850.n1900, inst_s15850.n1901, inst_s15850.n1902, inst_s15850.n1903, inst_s15850.n1904, inst_s15850.n1905, inst_s15850.n1906, inst_s15850.n1907, inst_s15850.n1908, inst_s15850.n1909, inst_s15850.n1910, inst_s15850.n1911, inst_s15850.n1912, inst_s15850.n1913, inst_s15850.n1914, inst_s15850.n1915, inst_s15850.n1916, inst_s15850.n1917, inst_s15850.n1918, inst_s15850.n1919, inst_s15850.n1920, inst_s15850.n1921, inst_s15850.n1922, inst_s15850.n1923, inst_s15850.n1924, inst_s15850.n1925, inst_s15850.n1926, inst_s15850.n1927, inst_s15850.n1928, inst_s15850.n1929, inst_s15850.n1930, inst_s15850.n1931, inst_s15850.n1932, inst_s15850.n1933, inst_s15850.n1934, inst_s15850.n1935, inst_s15850.n1936, inst_s15850.n1937, inst_s15850.n1938, inst_s15850.n1939, inst_s15850.n1940, inst_s15850.n1941, inst_s15850.n1942, inst_s15850.n1943, inst_s15850.n1944, inst_s15850.n1945, inst_s15850.n1946, inst_s15850.n1947, inst_s15850.n1948, inst_s15850.n1949, inst_s15850.n1950, inst_s15850.n1951, inst_s15850.n1952, inst_s15850.n1953, inst_s15850.n1954, inst_s15850.n1955, inst_s15850.n1956, inst_s15850.n1957, inst_s15850.n1958, inst_s15850.n1959, inst_s15850.n1960, inst_s15850.n1961, inst_s15850.n1962, inst_s15850.n1963, inst_s15850.n1964, inst_s15850.n1965, inst_s15850.n1966, inst_s15850.n1967, inst_s15850.n1968, inst_s15850.n1969, inst_s15850.n1970, inst_s15850.n1971, inst_s15850.n1972, inst_s15850.n1973, inst_s15850.n1974, inst_s15850.n1975, inst_s15850.n1976, inst_s15850.n1977, inst_s15850.n1978, inst_s15850.n1979, inst_s15850.n1980, inst_s15850.n1981, inst_s15850.n1982, inst_s15850.n1983, inst_s15850.n1984, inst_s15850.n1985, inst_s15850.n1986, inst_s15850.n1987, inst_s15850.n1988, inst_s15850.n3016, inst_s15850.n3017, inst_s15850.n3018, inst_s15850.n3019, inst_s15850.n3020, inst_s15850.n3022, inst_s15850.n3023, inst_s15850.n3024, inst_s15850.n3025, inst_s15850.n3026, inst_s15850.n3027, inst_s15850.n3029, inst_s15850.n3030, inst_s15850.n3031, inst_s15850.n3033, inst_s15850.n3034, inst_s15850.n3035, inst_s15850.n3036, inst_s15850.n3037, inst_s15850.n3038, inst_s15850.n3040, inst_s15850.n3041, inst_s15850.n3042, inst_s15850.n3044, inst_s15850.n3045, inst_s15850.n3046, inst_s15850.n3047, inst_s15850.n3048, inst_s15850.n3050, inst_s15850.n3051, inst_s15850.n3053, inst_s15850.n3054, inst_s15850.n3055, inst_s15850.n3056, inst_s15850.n3057, inst_s15850.n3058, inst_s15850.n3059, inst_s15850.n3061, inst_s15850.n3062, inst_s15850.n3064, inst_s15850.n3065, inst_s15850.Tg1, inst_s15850.Tg1_OUT1, inst_s15850.Tg1_OUT1234, inst_s15850.Tg1_OUT2, inst_s15850.Tg1_OUT3, inst_s15850.Tg1_OUT4, inst_s15850.Tg1_OUT5, inst_s15850.Tg1_OUT5678, inst_s15850.Tg1_OUT6, inst_s15850.Tg1_OUT7, inst_s15850.Tg1_OUT8, inst_s15850.Tg1_Trigger1, inst_s15850.Tg2, inst_s15850.Tg2_OUT1, inst_s15850.Tg2_OUT1234, inst_s15850.Tg2_OUT2, inst_s15850.Tg2_OUT3, inst_s15850.Tg2_OUT4, inst_s15850.Tg2_OUT5, inst_s15850.Tg2_OUT5678, inst_s15850.Tg2_OUT6, inst_s15850.Tg2_OUT7, inst_s15850.Tg2_OUT8, inst_s15850.Tg2_Trigger2, inst_s15850.Trigger_select);
        end
        $fclose(fptr);
        $finish;
    end
endmodule