`timescale 1ns / 1ps

`include "s38417_scan.v"

module tb_s38417;
    integer fptr;
    localparam Size = 1056768;
    reg [129:0] test_data [1056767:0];
    integer i = 0;

    reg CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;

    wire g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;

    `define in_data {g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se, test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9, test_si10, test_si11, test_si12, test_si13, test_si14, test_si15, test_si16, test_si17, test_si18, test_si19, test_si20, test_si21, test_si22, test_si23, test_si24, test_si25, test_si26, test_si27, test_si28, test_si29, test_si30, test_si31, test_si32, test_si33, test_si34, test_si35, test_si36, test_si37, test_si38, test_si39, test_si40, test_si41, test_si42, test_si43, test_si44, test_si45, test_si46, test_si47, test_si48, test_si49, test_si50, test_si51, test_si52, test_si53, test_si54, test_si55, test_si56, test_si57, test_si58, test_si59, test_si60, test_si61, test_si62, test_si63, test_si64, test_si65, test_si66, test_si67, test_si68, test_si69, test_si70, test_si71, test_si72, test_si73, test_si74, test_si75, test_si76, test_si77, test_si78, test_si79, test_si80, test_si81, test_si82, test_si83, test_si84, test_si85, test_si86, test_si87, test_si88, test_si89, test_si90, test_si91, test_si92, test_si93, test_si94, test_si95, test_si96, test_si97, test_si98, test_si99, test_si100}

    s38417 inst_s38417 (
    .CK (CK),
    .g1249 (g1249),
    .g1943 (g1943),
    .g2637 (g2637),
    .g3212 (g3212),
    .g3213 (g3213),
    .g3214 (g3214),
    .g3215 (g3215),
    .g3216 (g3216),
    .g3217 (g3217),
    .g3218 (g3218),
    .g3219 (g3219),
    .g3220 (g3220),
    .g3221 (g3221),
    .g3222 (g3222),
    .g3223 (g3223),
    .g3224 (g3224),
    .g3225 (g3225),
    .g3226 (g3226),
    .g3227 (g3227),
    .g3228 (g3228),
    .g3229 (g3229),
    .g3230 (g3230),
    .g3231 (g3231),
    .g3232 (g3232),
    .g3233 (g3233),
    .g3234 (g3234),
    .g51 (g51),
    .g563 (g563),
    .test_se (test_se),
    .test_si1 (test_si1),
    .test_si2 (test_si2),
    .test_si3 (test_si3),
    .test_si4 (test_si4),
    .test_si5 (test_si5),
    .test_si6 (test_si6),
    .test_si7 (test_si7),
    .test_si8 (test_si8),
    .test_si9 (test_si9),
    .test_si10 (test_si10),
    .test_si11 (test_si11),
    .test_si12 (test_si12),
    .test_si13 (test_si13),
    .test_si14 (test_si14),
    .test_si15 (test_si15),
    .test_si16 (test_si16),
    .test_si17 (test_si17),
    .test_si18 (test_si18),
    .test_si19 (test_si19),
    .test_si20 (test_si20),
    .test_si21 (test_si21),
    .test_si22 (test_si22),
    .test_si23 (test_si23),
    .test_si24 (test_si24),
    .test_si25 (test_si25),
    .test_si26 (test_si26),
    .test_si27 (test_si27),
    .test_si28 (test_si28),
    .test_si29 (test_si29),
    .test_si30 (test_si30),
    .test_si31 (test_si31),
    .test_si32 (test_si32),
    .test_si33 (test_si33),
    .test_si34 (test_si34),
    .test_si35 (test_si35),
    .test_si36 (test_si36),
    .test_si37 (test_si37),
    .test_si38 (test_si38),
    .test_si39 (test_si39),
    .test_si40 (test_si40),
    .test_si41 (test_si41),
    .test_si42 (test_si42),
    .test_si43 (test_si43),
    .test_si44 (test_si44),
    .test_si45 (test_si45),
    .test_si46 (test_si46),
    .test_si47 (test_si47),
    .test_si48 (test_si48),
    .test_si49 (test_si49),
    .test_si50 (test_si50),
    .test_si51 (test_si51),
    .test_si52 (test_si52),
    .test_si53 (test_si53),
    .test_si54 (test_si54),
    .test_si55 (test_si55),
    .test_si56 (test_si56),
    .test_si57 (test_si57),
    .test_si58 (test_si58),
    .test_si59 (test_si59),
    .test_si60 (test_si60),
    .test_si61 (test_si61),
    .test_si62 (test_si62),
    .test_si63 (test_si63),
    .test_si64 (test_si64),
    .test_si65 (test_si65),
    .test_si66 (test_si66),
    .test_si67 (test_si67),
    .test_si68 (test_si68),
    .test_si69 (test_si69),
    .test_si70 (test_si70),
    .test_si71 (test_si71),
    .test_si72 (test_si72),
    .test_si73 (test_si73),
    .test_si74 (test_si74),
    .test_si75 (test_si75),
    .test_si76 (test_si76),
    .test_si77 (test_si77),
    .test_si78 (test_si78),
    .test_si79 (test_si79),
    .test_si80 (test_si80),
    .test_si81 (test_si81),
    .test_si82 (test_si82),
    .test_si83 (test_si83),
    .test_si84 (test_si84),
    .test_si85 (test_si85),
    .test_si86 (test_si86),
    .test_si87 (test_si87),
    .test_si88 (test_si88),
    .test_si89 (test_si89),
    .test_si90 (test_si90),
    .test_si91 (test_si91),
    .test_si92 (test_si92),
    .test_si93 (test_si93),
    .test_si94 (test_si94),
    .test_si95 (test_si95),
    .test_si96 (test_si96),
    .test_si97 (test_si97),
    .test_si98 (test_si98),
    .test_si99 (test_si99),
    .test_si100 (test_si100));


    initial begin
    // $dumpfile("s15850.vcd");
    // $dumpvars(0, tb_s15850);
    fptr = $fopen("data_out.txt", "w");

    $readmemb("s38417_4096samples.vec", test_data);
    for (i=0; i<Size; i = i + 1) begin
        `in_data = test_data[i]; #10;

        $fwrite(fptr, "%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d%d\n", inst_s38417.N690, inst_s38417.N995, inst_s38417.g2950, inst_s38417.g2883, inst_s38417.g2888, inst_s38417.g2896, inst_s38417.g2892, inst_s38417.g2903, inst_s38417.g2900, inst_s38417.g2908, inst_s38417.g2912, inst_s38417.g2917, inst_s38417.g2924, inst_s38417.g2920, inst_s38417.g2879, inst_s38417.g2934, inst_s38417.g2935, inst_s38417.g2938, inst_s38417.g2941, inst_s38417.g2944, inst_s38417.g2947, inst_s38417.g2953, inst_s38417.g2956, inst_s38417.g2959, inst_s38417.g2962, inst_s38417.g2963, inst_s38417.g2969, inst_s38417.g2972, inst_s38417.g2975, inst_s38417.g2978, inst_s38417.g2981, inst_s38417.g2874, inst_s38417.g1506, inst_s38417.g1501, inst_s38417.g1496, inst_s38417.g1491, inst_s38417.g1486, inst_s38417.g1481, inst_s38417.g1476, inst_s38417.g1471, inst_s38417.g2877, inst_s38417.g8251, inst_s38417.g813, inst_s38417.g809, inst_s38417.g805, inst_s38417.g801, inst_s38417.g797, inst_s38417.g793, inst_s38417.g789, inst_s38417.g785, inst_s38417.g7519, inst_s38417.g2873, inst_s38417.g125, inst_s38417.g121, inst_s38417.g117, inst_s38417.g113, inst_s38417.g109, inst_s38417.g105, inst_s38417.g101, inst_s38417.g4450, inst_s38417.g97, inst_s38417.g2857, inst_s38417.g2200, inst_s38417.g2195, inst_s38417.g2190, inst_s38417.g2185, inst_s38417.g2180, inst_s38417.g2175, inst_s38417.g2170, inst_s38417.g2165, inst_s38417.g2878, inst_s38417.g3129, inst_s38417.g3117, inst_s38417.g3109, inst_s38417.g3211, inst_s38417.g3084, inst_s38417.g3085, inst_s38417.g3086, inst_s38417.g3087, inst_s38417.g3091, inst_s38417.g3092, inst_s38417.g3093, inst_s38417.g3094, inst_s38417.g3095, inst_s38417.g3096, inst_s38417.g3097, inst_s38417.g3098, inst_s38417.g3099, inst_s38417.g3100, inst_s38417.g3102, inst_s38417.g3103, inst_s38417.g3104, inst_s38417.g3105, inst_s38417.g3106, inst_s38417.g3107, inst_s38417.g3108, inst_s38417.g3155, inst_s38417.g3158, inst_s38417.g3161, inst_s38417.g3164, inst_s38417.g3167, inst_s38417.g3170, inst_s38417.g3173, inst_s38417.g3176, inst_s38417.g3182, inst_s38417.g3185, inst_s38417.g3088, inst_s38417.g3197, inst_s38417.g3201, inst_s38417.g3204, inst_s38417.g3207, inst_s38417.g3188, inst_s38417.g3133, inst_s38417.g3128, inst_s38417.g3124, inst_s38417.g3112, inst_s38417.g3110, inst_s38417.g3111, inst_s38417.g3151, inst_s38417.g3142, inst_s38417.g185, inst_s38417.g138, inst_s38417.g165, inst_s38417.g130, inst_s38417.g131, inst_s38417.g129, inst_s38417.g133, inst_s38417.g134, inst_s38417.g132, inst_s38417.g142, inst_s38417.g143, inst_s38417.g141, inst_s38417.g145, inst_s38417.g146, inst_s38417.g148, inst_s38417.g149, inst_s38417.g147, inst_s38417.g151, inst_s38417.g152, inst_s38417.g150, inst_s38417.g154, inst_s38417.g155, inst_s38417.g153, inst_s38417.g157, inst_s38417.g158, inst_s38417.g156, inst_s38417.g160, inst_s38417.g161, inst_s38417.g159, inst_s38417.g164, inst_s38417.g162, inst_s38417.g169, inst_s38417.g170, inst_s38417.g168, inst_s38417.g172, inst_s38417.g173, inst_s38417.g171, inst_s38417.g175, inst_s38417.g176, inst_s38417.g174, inst_s38417.g178, inst_s38417.g179, inst_s38417.g177, inst_s38417.g186, inst_s38417.g192, inst_s38417.g231, inst_s38417.g234, inst_s38417.g237, inst_s38417.g195, inst_s38417.g198, inst_s38417.g201, inst_s38417.g240, inst_s38417.g243, inst_s38417.g246, inst_s38417.g204, inst_s38417.g207, inst_s38417.g210, inst_s38417.g249, inst_s38417.g252, inst_s38417.g213, inst_s38417.g216, inst_s38417.g219, inst_s38417.g258, inst_s38417.g261, inst_s38417.g264, inst_s38417.g222, inst_s38417.g225, inst_s38417.g228, inst_s38417.g267, inst_s38417.g270, inst_s38417.g273, inst_s38417.g92, inst_s38417.g88, inst_s38417.g83, inst_s38417.g74, inst_s38417.g70, inst_s38417.g65, inst_s38417.g61, inst_s38417.g56, inst_s38417.g52, inst_s38417.g180, inst_s38417.g181, inst_s38417.g276, inst_s38417.g401, inst_s38417.g309, inst_s38417.g354, inst_s38417.g343, inst_s38417.g369, inst_s38417.g358, inst_s38417.g361, inst_s38417.g384, inst_s38417.g373, inst_s38417.g376, inst_s38417.g398, inst_s38417.g388, inst_s38417.g391, inst_s38417.g408, inst_s38417.g411, inst_s38417.g414, inst_s38417.g417, inst_s38417.g420, inst_s38417.g423, inst_s38417.g428, inst_s38417.g426, inst_s38417.g429, inst_s38417.g432, inst_s38417.g435, inst_s38417.g438, inst_s38417.g441, inst_s38417.g444, inst_s38417.g448, inst_s38417.g449, inst_s38417.g447, inst_s38417.g312, inst_s38417.g313, inst_s38417.g314, inst_s38417.g315, inst_s38417.g317, inst_s38417.g318, inst_s38417.g319, inst_s38417.g320, inst_s38417.g322, inst_s38417.g323, inst_s38417.g321, inst_s38417.g403, inst_s38417.g404, inst_s38417.g402, inst_s38417.g450, inst_s38417.g452, inst_s38417.g454, inst_s38417.g280, inst_s38417.g282, inst_s38417.g284, inst_s38417.g286, inst_s38417.g288, inst_s38417.g290, inst_s38417.g305, inst_s38417.g349, inst_s38417.g350, inst_s38417.g351, inst_s38417.g352, inst_s38417.g353, inst_s38417.g357, inst_s38417.g364, inst_s38417.g365, inst_s38417.g366, inst_s38417.g367, inst_s38417.g368, inst_s38417.g372, inst_s38417.g379, inst_s38417.g380, inst_s38417.g381, inst_s38417.g383, inst_s38417.g387, inst_s38417.g394, inst_s38417.g395, inst_s38417.g396, inst_s38417.g397, inst_s38417.g324, inst_s38417.g337, inst_s38417.g545, inst_s38417.g551, inst_s38417.g550, inst_s38417.g554, inst_s38417.g557, inst_s38417.g513, inst_s38417.g523, inst_s38417.g524, inst_s38417.g564, inst_s38417.g569, inst_s38417.g570, inst_s38417.g571, inst_s38417.g572, inst_s38417.g573, inst_s38417.g574, inst_s38417.g565, inst_s38417.g566, inst_s38417.g567, inst_s38417.g568, inst_s38417.g489, inst_s38417.g7909, inst_s38417.g485, inst_s38417.g486, inst_s38417.g487, inst_s38417.g488, inst_s38417.g455, inst_s38417.g458, inst_s38417.g461, inst_s38417.g477, inst_s38417.g478, inst_s38417.g479, inst_s38417.g480, inst_s38417.g484, inst_s38417.g464, inst_s38417.g465, inst_s38417.g471, inst_s38417.g528, inst_s38417.g535, inst_s38417.g542, inst_s38417.g543, inst_s38417.g544, inst_s38417.g548, inst_s38417.g549, inst_s38417.g499, inst_s38417.g558, inst_s38417.g559, inst_s38417.g576, inst_s38417.g577, inst_s38417.g575, inst_s38417.g579, inst_s38417.g578, inst_s38417.g582, inst_s38417.g583, inst_s38417.g581, inst_s38417.g585, inst_s38417.g586, inst_s38417.g584, inst_s38417.g587, inst_s38417.g590, inst_s38417.g593, inst_s38417.g596, inst_s38417.g599, inst_s38417.g602, inst_s38417.g614, inst_s38417.g617, inst_s38417.g605, inst_s38417.g608, inst_s38417.g611, inst_s38417.g490, inst_s38417.g493, inst_s38417.g496, inst_s38417.g506, inst_s38417.g525, inst_s38417.g536, inst_s38417.g537, inst_s38417.g538, inst_s38417.g629, inst_s38417.g630, inst_s38417.g659, inst_s38417.g640, inst_s38417.g633, inst_s38417.g653, inst_s38417.g646, inst_s38417.g660, inst_s38417.g672, inst_s38417.g679, inst_s38417.g686, inst_s38417.g692, inst_s38417.g699, inst_s38417.g700, inst_s38417.g698, inst_s38417.g702, inst_s38417.g703, inst_s38417.g701, inst_s38417.g705, inst_s38417.g706, inst_s38417.g704, inst_s38417.g708, inst_s38417.g709, inst_s38417.g707, inst_s38417.g712, inst_s38417.g710, inst_s38417.g714, inst_s38417.g715, inst_s38417.g713, inst_s38417.g717, inst_s38417.g718, inst_s38417.g716, inst_s38417.g720, inst_s38417.g721, inst_s38417.g719, inst_s38417.g723, inst_s38417.g724, inst_s38417.g722, inst_s38417.g726, inst_s38417.g725, inst_s38417.g729, inst_s38417.g730, inst_s38417.g728, inst_s38417.g732, inst_s38417.g733, inst_s38417.g731, inst_s38417.g735, inst_s38417.g736, inst_s38417.g734, inst_s38417.g738, inst_s38417.g739, inst_s38417.g737, inst_s38417.g818, inst_s38417.g819, inst_s38417.g817, inst_s38417.g821, inst_s38417.g822, inst_s38417.g820, inst_s38417.g830, inst_s38417.g831, inst_s38417.g829, inst_s38417.g833, inst_s38417.g834, inst_s38417.g832, inst_s38417.g836, inst_s38417.g837, inst_s38417.g835, inst_s38417.g840, inst_s38417.g838, inst_s38417.g842, inst_s38417.g843, inst_s38417.g841, inst_s38417.g845, inst_s38417.g846, inst_s38417.g844, inst_s38417.g848, inst_s38417.g849, inst_s38417.g847, inst_s38417.g851, inst_s38417.g852, inst_s38417.g850, inst_s38417.g857, inst_s38417.g856, inst_s38417.g860, inst_s38417.g861, inst_s38417.g859, inst_s38417.g863, inst_s38417.g864, inst_s38417.g862, inst_s38417.g866, inst_s38417.g867, inst_s38417.g865, inst_s38417.g873, inst_s38417.g876, inst_s38417.g879, inst_s38417.g918, inst_s38417.g921, inst_s38417.g882, inst_s38417.g885, inst_s38417.g888, inst_s38417.g927, inst_s38417.g930, inst_s38417.g933, inst_s38417.g891, inst_s38417.g894, inst_s38417.g897, inst_s38417.g936, inst_s38417.g939, inst_s38417.g942, inst_s38417.g900, inst_s38417.g903, inst_s38417.g906, inst_s38417.g948, inst_s38417.g951, inst_s38417.g909, inst_s38417.g912, inst_s38417.g915, inst_s38417.g954, inst_s38417.g957, inst_s38417.g960, inst_s38417.g780, inst_s38417.g776, inst_s38417.g771, inst_s38417.g767, inst_s38417.g762, inst_s38417.g758, inst_s38417.g753, inst_s38417.g744, inst_s38417.g740, inst_s38417.g868, inst_s38417.g869, inst_s38417.g963, inst_s38417.g1092, inst_s38417.g1088, inst_s38417.g996, inst_s38417.g1041, inst_s38417.g1030, inst_s38417.g1033, inst_s38417.g1056, inst_s38417.g1045, inst_s38417.g1048, inst_s38417.g1060, inst_s38417.g1063, inst_s38417.g1085, inst_s38417.g1075, inst_s38417.g1078, inst_s38417.g1095, inst_s38417.g1098, inst_s38417.g1101, inst_s38417.g1104, inst_s38417.g1107, inst_s38417.g1110, inst_s38417.g1114, inst_s38417.g1115, inst_s38417.g1113, inst_s38417.g1116, inst_s38417.g1122, inst_s38417.g1125, inst_s38417.g1128, inst_s38417.g1131, inst_s38417.g1135, inst_s38417.g1136, inst_s38417.g1134, inst_s38417.g999, inst_s38417.g1000, inst_s38417.g1001, inst_s38417.g1002, inst_s38417.g1003, inst_s38417.g1004, inst_s38417.g1005, inst_s38417.g1006, inst_s38417.g1009, inst_s38417.g1010, inst_s38417.g1008, inst_s38417.g1090, inst_s38417.g1091, inst_s38417.g1089, inst_s38417.g1137, inst_s38417.g1139, inst_s38417.g1141, inst_s38417.g967, inst_s38417.g969, inst_s38417.g971, inst_s38417.g973, inst_s38417.g975, inst_s38417.g977, inst_s38417.g986, inst_s38417.g992, inst_s38417.g1029, inst_s38417.g1036, inst_s38417.g1037, inst_s38417.g1038, inst_s38417.g1040, inst_s38417.g1044, inst_s38417.g1051, inst_s38417.g1052, inst_s38417.g1053, inst_s38417.g1054, inst_s38417.g1055, inst_s38417.g1059, inst_s38417.g1066, inst_s38417.g1067, inst_s38417.g1068, inst_s38417.g1069, inst_s38417.g1070, inst_s38417.g1074, inst_s38417.g1081, inst_s38417.g1083, inst_s38417.g1084, inst_s38417.g1011, inst_s38417.g1024, inst_s38417.g1231, inst_s38417.g1237, inst_s38417.g1236, inst_s38417.g1240, inst_s38417.g1243, inst_s38417.g1196, inst_s38417.g1199, inst_s38417.g1209, inst_s38417.g1210, inst_s38417.g1255, inst_s38417.g1256, inst_s38417.g1257, inst_s38417.g1258, inst_s38417.g1259, inst_s38417.g1260, inst_s38417.g1251, inst_s38417.g1252, inst_s38417.g1253, inst_s38417.g1254, inst_s38417.g1176, inst_s38417.g1172, inst_s38417.g1173, inst_s38417.g1175, inst_s38417.g1142, inst_s38417.g1145, inst_s38417.g1148, inst_s38417.g1164, inst_s38417.g1165, inst_s38417.g1166, inst_s38417.g1167, inst_s38417.g1171, inst_s38417.g1151, inst_s38417.g1152, inst_s38417.g1155, inst_s38417.g1158, inst_s38417.g1214, inst_s38417.g1221, inst_s38417.g1229, inst_s38417.g1235, inst_s38417.g1186, inst_s38417.g1244, inst_s38417.g1245, inst_s38417.g1262, inst_s38417.g1263, inst_s38417.g1261, inst_s38417.g1265, inst_s38417.g1266, inst_s38417.g1264, inst_s38417.g1268, inst_s38417.g1269, inst_s38417.g1271, inst_s38417.g1272, inst_s38417.g1270, inst_s38417.g1273, inst_s38417.g1276, inst_s38417.g1279, inst_s38417.g1282, inst_s38417.g1285, inst_s38417.g1288, inst_s38417.g1300, inst_s38417.g1303, inst_s38417.g1306, inst_s38417.g1291, inst_s38417.g1294, inst_s38417.g1297, inst_s38417.g1180, inst_s38417.g1183, inst_s38417.g1192, inst_s38417.g1211, inst_s38417.g1222, inst_s38417.g1223, inst_s38417.g1224, inst_s38417.g1315, inst_s38417.g1316, inst_s38417.g1345, inst_s38417.g1326, inst_s38417.g1319, inst_s38417.g1339, inst_s38417.g1332, inst_s38417.g1346, inst_s38417.g1358, inst_s38417.g1352, inst_s38417.g1365, inst_s38417.g1372, inst_s38417.g1378, inst_s38417.g1386, inst_s38417.g1384, inst_s38417.g1388, inst_s38417.g1389, inst_s38417.g1387, inst_s38417.g1391, inst_s38417.g1392, inst_s38417.g1390, inst_s38417.g1394, inst_s38417.g1395, inst_s38417.g1393, inst_s38417.g1397, inst_s38417.g1398, inst_s38417.g1396, inst_s38417.g1400, inst_s38417.g1399, inst_s38417.g1403, inst_s38417.g1404, inst_s38417.g1402, inst_s38417.g1406, inst_s38417.g1407, inst_s38417.g1405, inst_s38417.g1409, inst_s38417.g1410, inst_s38417.g1408, inst_s38417.g1412, inst_s38417.g1413, inst_s38417.g1411, inst_s38417.g1415, inst_s38417.g1416, inst_s38417.g1418, inst_s38417.g1419, inst_s38417.g1417, inst_s38417.g1421, inst_s38417.g1422, inst_s38417.g1420, inst_s38417.g1424, inst_s38417.g1425, inst_s38417.g1423, inst_s38417.g1520, inst_s38417.g1547, inst_s38417.g1512, inst_s38417.g1513, inst_s38417.g1511, inst_s38417.g1516, inst_s38417.g1514, inst_s38417.g1524, inst_s38417.g1525, inst_s38417.g1523, inst_s38417.g1527, inst_s38417.g1528, inst_s38417.g1526, inst_s38417.g1530, inst_s38417.g1531, inst_s38417.g1529, inst_s38417.g1533, inst_s38417.g1534, inst_s38417.g1532, inst_s38417.g1536, inst_s38417.g1535, inst_s38417.g1539, inst_s38417.g1540, inst_s38417.g1538, inst_s38417.g1542, inst_s38417.g1543, inst_s38417.g1541, inst_s38417.g1545, inst_s38417.g1546, inst_s38417.g1544, inst_s38417.g1551, inst_s38417.g1552, inst_s38417.g1550, inst_s38417.g1554, inst_s38417.g1555, inst_s38417.g1557, inst_s38417.g1558, inst_s38417.g1556, inst_s38417.g1560, inst_s38417.g1561, inst_s38417.g1559, inst_s38417.g1567, inst_s38417.g1570, inst_s38417.g1573, inst_s38417.g1612, inst_s38417.g1615, inst_s38417.g1618, inst_s38417.g1576, inst_s38417.g1579, inst_s38417.g1582, inst_s38417.g1624, inst_s38417.g1627, inst_s38417.g1585, inst_s38417.g1588, inst_s38417.g1591, inst_s38417.g1630, inst_s38417.g1633, inst_s38417.g1636, inst_s38417.g1594, inst_s38417.g1597, inst_s38417.g1600, inst_s38417.g1639, inst_s38417.g1642, inst_s38417.g1645, inst_s38417.g1603, inst_s38417.g1609, inst_s38417.g1648, inst_s38417.g1651, inst_s38417.g1654, inst_s38417.g1466, inst_s38417.g1462, inst_s38417.g1457, inst_s38417.g1453, inst_s38417.g1448, inst_s38417.g1444, inst_s38417.g1439, inst_s38417.g1435, inst_s38417.g1430, inst_s38417.g1426, inst_s38417.g1562, inst_s38417.g5612, inst_s38417.g1563, inst_s38417.g1657, inst_s38417.g1786, inst_s38417.g1782, inst_s38417.g1690, inst_s38417.g1735, inst_s38417.g1724, inst_s38417.g1727, inst_s38417.g1750, inst_s38417.g1739, inst_s38417.g1742, inst_s38417.g1765, inst_s38417.g1754, inst_s38417.g1757, inst_s38417.g1779, inst_s38417.g1772, inst_s38417.g1789, inst_s38417.g1792, inst_s38417.g1795, inst_s38417.g1798, inst_s38417.g1801, inst_s38417.g1804, inst_s38417.g1808, inst_s38417.g1809, inst_s38417.g1807, inst_s38417.g1810, inst_s38417.g1813, inst_s38417.g1816, inst_s38417.g1819, inst_s38417.g1822, inst_s38417.g1829, inst_s38417.g1830, inst_s38417.g1828, inst_s38417.g1693, inst_s38417.g1694, inst_s38417.g1695, inst_s38417.g1696, inst_s38417.g1697, inst_s38417.g1698, inst_s38417.g1699, inst_s38417.g1700, inst_s38417.g1701, inst_s38417.g1703, inst_s38417.g1704, inst_s38417.g1702, inst_s38417.g1785, inst_s38417.g1783, inst_s38417.g1831, inst_s38417.g1833, inst_s38417.g1835, inst_s38417.g1661, inst_s38417.g1663, inst_s38417.g1665, inst_s38417.g1667, inst_s38417.g1669, inst_s38417.g1671, inst_s38417.g1680, inst_s38417.g1686, inst_s38417.g1723, inst_s38417.g1730, inst_s38417.g1731, inst_s38417.g1732, inst_s38417.g1733, inst_s38417.g1734, inst_s38417.g1738, inst_s38417.g1745, inst_s38417.g1747, inst_s38417.g1748, inst_s38417.g1749, inst_s38417.g1753, inst_s38417.g1760, inst_s38417.g1761, inst_s38417.g1762, inst_s38417.g1763, inst_s38417.g1764, inst_s38417.g1768, inst_s38417.g1775, inst_s38417.g1776, inst_s38417.g1777, inst_s38417.g1778, inst_s38417.g1705, inst_s38417.g5695, inst_s38417.g1718, inst_s38417.g1925, inst_s38417.g1931, inst_s38417.g1930, inst_s38417.g1934, inst_s38417.g1937, inst_s38417.g1890, inst_s38417.g1893, inst_s38417.g1903, inst_s38417.g1904, inst_s38417.g1944, inst_s38417.g1949, inst_s38417.g1950, inst_s38417.g1951, inst_s38417.g1953, inst_s38417.g1954, inst_s38417.g1945, inst_s38417.g1946, inst_s38417.g1947, inst_s38417.g1948, inst_s38417.g1870, inst_s38417.g1866, inst_s38417.g1867, inst_s38417.g1868, inst_s38417.g1869, inst_s38417.g1836, inst_s38417.g1842, inst_s38417.g1858, inst_s38417.g1859, inst_s38417.g1860, inst_s38417.g1861, inst_s38417.g1865, inst_s38417.g1845, inst_s38417.g1846, inst_s38417.g1849, inst_s38417.g1852, inst_s38417.g1908, inst_s38417.g1915, inst_s38417.g1922, inst_s38417.g1923, inst_s38417.g1929, inst_s38417.g1880, inst_s38417.g1938, inst_s38417.g1939, inst_s38417.g1956, inst_s38417.g1957, inst_s38417.g1955, inst_s38417.g1959, inst_s38417.g1960, inst_s38417.g1958, inst_s38417.g1962, inst_s38417.g1963, inst_s38417.g1961, inst_s38417.g1966, inst_s38417.g1964, inst_s38417.g1967, inst_s38417.g1970, inst_s38417.g1973, inst_s38417.g1976, inst_s38417.g1979, inst_s38417.g1982, inst_s38417.g1994, inst_s38417.g1997, inst_s38417.g2000, inst_s38417.g1985, inst_s38417.g1988, inst_s38417.g1991, inst_s38417.g1874, inst_s38417.g1877, inst_s38417.g1886, inst_s38417.g1905, inst_s38417.g1916, inst_s38417.g1917, inst_s38417.g2009, inst_s38417.g2010, inst_s38417.g2039, inst_s38417.g2020, inst_s38417.g2013, inst_s38417.g2033, inst_s38417.g2026, inst_s38417.g2040, inst_s38417.g2052, inst_s38417.g2046, inst_s38417.g2059, inst_s38417.g2072, inst_s38417.g2079, inst_s38417.g2080, inst_s38417.g2078, inst_s38417.g2082, inst_s38417.g2083, inst_s38417.g2081, inst_s38417.g2085, inst_s38417.g2086, inst_s38417.g2084, inst_s38417.g2088, inst_s38417.g2089, inst_s38417.g2087, inst_s38417.g2091, inst_s38417.g2090, inst_s38417.g2094, inst_s38417.g2095, inst_s38417.g2093, inst_s38417.g2097, inst_s38417.g2098, inst_s38417.g2096, inst_s38417.g2100, inst_s38417.g2101, inst_s38417.g2099, inst_s38417.g2103, inst_s38417.g2104, inst_s38417.g2102, inst_s38417.g2106, inst_s38417.g2105, inst_s38417.g2109, inst_s38417.g2110, inst_s38417.g2108, inst_s38417.g2112, inst_s38417.g2113, inst_s38417.g2111, inst_s38417.g2115, inst_s38417.g2116, inst_s38417.g2114, inst_s38417.g2118, inst_s38417.g2119, inst_s38417.g2117, inst_s38417.g2214, inst_s38417.g7084, inst_s38417.g2241, inst_s38417.g2206, inst_s38417.g2207, inst_s38417.g2205, inst_s38417.g2209, inst_s38417.g2210, inst_s38417.g2208, inst_s38417.g2218, inst_s38417.g2219, inst_s38417.g2217, inst_s38417.g2221, inst_s38417.g2222, inst_s38417.g2220, inst_s38417.g2224, inst_s38417.g2223, inst_s38417.g2227, inst_s38417.g2228, inst_s38417.g2226, inst_s38417.g2230, inst_s38417.g2231, inst_s38417.g2229, inst_s38417.g2233, inst_s38417.g2234, inst_s38417.g2232, inst_s38417.g2236, inst_s38417.g2237, inst_s38417.g2235, inst_s38417.g2239, inst_s38417.g2238, inst_s38417.g2245, inst_s38417.g2246, inst_s38417.g2244, inst_s38417.g2248, inst_s38417.g2249, inst_s38417.g2247, inst_s38417.g2251, inst_s38417.g2252, inst_s38417.g2250, inst_s38417.g2254, inst_s38417.g2255, inst_s38417.g2253, inst_s38417.g2261, inst_s38417.g2267, inst_s38417.g2306, inst_s38417.g2309, inst_s38417.g2312, inst_s38417.g2270, inst_s38417.g2273, inst_s38417.g2276, inst_s38417.g2315, inst_s38417.g2318, inst_s38417.g2321, inst_s38417.g2279, inst_s38417.g2282, inst_s38417.g2285, inst_s38417.g2324, inst_s38417.g2330, inst_s38417.g2288, inst_s38417.g2291, inst_s38417.g2294, inst_s38417.g2333, inst_s38417.g2336, inst_s38417.g2339, inst_s38417.g2297, inst_s38417.g2300, inst_s38417.g2303, inst_s38417.g2342, inst_s38417.g2345, inst_s38417.g2348, inst_s38417.g2160, inst_s38417.g2151, inst_s38417.g2147, inst_s38417.g2142, inst_s38417.g2138, inst_s38417.g2133, inst_s38417.g2129, inst_s38417.g2124, inst_s38417.g2120, inst_s38417.g2256, inst_s38417.g2257, inst_s38417.g2351, inst_s38417.g2480, inst_s38417.g2476, inst_s38417.g2429, inst_s38417.g2418, inst_s38417.g2421, inst_s38417.g2444, inst_s38417.g2433, inst_s38417.g2436, inst_s38417.g2459, inst_s38417.g2448, inst_s38417.g2451, inst_s38417.g2473, inst_s38417.g2463, inst_s38417.g2466, inst_s38417.g2483, inst_s38417.g2486, inst_s38417.g2492, inst_s38417.g2495, inst_s38417.g2498, inst_s38417.g2502, inst_s38417.g2503, inst_s38417.g2501, inst_s38417.g2504, inst_s38417.g2507, inst_s38417.g2510, inst_s38417.g2513, inst_s38417.g2516, inst_s38417.g2519, inst_s38417.g2523, inst_s38417.g2524, inst_s38417.g2387, inst_s38417.g2388, inst_s38417.g2389, inst_s38417.g2390, inst_s38417.g2391, inst_s38417.g2392, inst_s38417.g2393, inst_s38417.g2394, inst_s38417.g2395, inst_s38417.g2397, inst_s38417.g2398, inst_s38417.g2396, inst_s38417.g2478, inst_s38417.g2479, inst_s38417.g2525, inst_s38417.g2527, inst_s38417.g2529, inst_s38417.g2355, inst_s38417.g2357, inst_s38417.g2359, inst_s38417.g2361, inst_s38417.g2365, inst_s38417.g2374, inst_s38417.g2380, inst_s38417.g2417, inst_s38417.g2424, inst_s38417.g2425, inst_s38417.g2426, inst_s38417.g2427, inst_s38417.g2428, inst_s38417.g2432, inst_s38417.g2439, inst_s38417.g2441, inst_s38417.g2442, inst_s38417.g2443, inst_s38417.g2447, inst_s38417.g2454, inst_s38417.g2455, inst_s38417.g2456, inst_s38417.g2457, inst_s38417.g2458, inst_s38417.g2462, inst_s38417.g2469, inst_s38417.g2470, inst_s38417.g2471, inst_s38417.g2472, inst_s38417.g2412, inst_s38417.g2619, inst_s38417.g2625, inst_s38417.g2624, inst_s38417.g2628, inst_s38417.g2631, inst_s38417.g2584, inst_s38417.g2587, inst_s38417.g2597, inst_s38417.g2598, inst_s38417.g2638, inst_s38417.g2643, inst_s38417.g2645, inst_s38417.g2646, inst_s38417.g2647, inst_s38417.g2648, inst_s38417.g2639, inst_s38417.g2640, inst_s38417.g2641, inst_s38417.g2642, inst_s38417.g2564, inst_s38417.g2560, inst_s38417.g2561, inst_s38417.g2562, inst_s38417.g2530, inst_s38417.g2533, inst_s38417.g2536, inst_s38417.g2552, inst_s38417.g2553, inst_s38417.g2554, inst_s38417.g2555, inst_s38417.g2559, inst_s38417.g2539, inst_s38417.g2540, inst_s38417.g2543, inst_s38417.g2546, inst_s38417.g2602, inst_s38417.g2609, inst_s38417.g2617, inst_s38417.g2623, inst_s38417.g2574, inst_s38417.g2632, inst_s38417.g2633, inst_s38417.g2650, inst_s38417.g2651, inst_s38417.g2649, inst_s38417.g2653, inst_s38417.g2654, inst_s38417.g2652, inst_s38417.g2656, inst_s38417.g2655, inst_s38417.g2659, inst_s38417.g2660, inst_s38417.g2658, inst_s38417.g2661, inst_s38417.g2664, inst_s38417.g2667, inst_s38417.g2670, inst_s38417.g2673, inst_s38417.g2676, inst_s38417.g2688, inst_s38417.g2691, inst_s38417.g2694, inst_s38417.g2679, inst_s38417.g2685, inst_s38417.g2565, inst_s38417.g2568, inst_s38417.g2571, inst_s38417.g2580, inst_s38417.g2599, inst_s38417.g2611, inst_s38417.g2612, inst_s38417.g2703, inst_s38417.g2704, inst_s38417.g2733, inst_s38417.g2714, inst_s38417.g2707, inst_s38417.g2727, inst_s38417.g2720, inst_s38417.g2734, inst_s38417.g2746, inst_s38417.g2753, inst_s38417.g2760, inst_s38417.g2766, inst_s38417.g2773, inst_s38417.g2774, inst_s38417.g2772, inst_s38417.g2776, inst_s38417.g2777, inst_s38417.g2775, inst_s38417.g2779, inst_s38417.g2780, inst_s38417.g2778, inst_s38417.g2782, inst_s38417.g2783, inst_s38417.g2785, inst_s38417.g2786, inst_s38417.g2784, inst_s38417.g2788, inst_s38417.g2789, inst_s38417.g2787, inst_s38417.g2791, inst_s38417.g2792, inst_s38417.g2790, inst_s38417.g2794, inst_s38417.g2795, inst_s38417.g2793, inst_s38417.g2797, inst_s38417.g2798, inst_s38417.g2800, inst_s38417.g2801, inst_s38417.g2799, inst_s38417.g2803, inst_s38417.g2804, inst_s38417.g2802, inst_s38417.g2806, inst_s38417.g2807, inst_s38417.g2805, inst_s38417.g2809, inst_s38417.g2810, inst_s38417.g2808, inst_s38417.g2812, inst_s38417.g2813, inst_s38417.g3080, inst_s38417.g3043, inst_s38417.g3044, inst_s38417.g3045, inst_s38417.g3046, inst_s38417.g3047, inst_s38417.g3048, inst_s38417.g3049, inst_s38417.g3050, inst_s38417.g3051, inst_s38417.g3052, inst_s38417.g3053, inst_s38417.g3056, inst_s38417.g3057, inst_s38417.g3058, inst_s38417.g3059, inst_s38417.g3060, inst_s38417.g3061, inst_s38417.g3062, inst_s38417.g3063, inst_s38417.g3064, inst_s38417.g3065, inst_s38417.g3066, inst_s38417.g3067, inst_s38417.g3068, inst_s38417.g3069, inst_s38417.g3071, inst_s38417.g3072, inst_s38417.g3073, inst_s38417.g3074, inst_s38417.g3075, inst_s38417.g3076, inst_s38417.g3077, inst_s38417.g3078, inst_s38417.g2997, inst_s38417.g2993, inst_s38417.g3006, inst_s38417.g3002, inst_s38417.g3013, inst_s38417.g3024, inst_s38417.g3018, inst_s38417.g3028, inst_s38417.g3036, inst_s38417.g3032, inst_s38417.g2987, inst_s38417.g8270, inst_s38417.g3083, inst_s38417.g2990, inst_s38417.g8258, inst_s38417.g13149, inst_s38417.g13111, inst_s38417.g13155, inst_s38417.g13160, inst_s38417.g13124, inst_s38417.g13164, inst_s38417.g12487, inst_s38417.g13171, inst_s38417.g13135, inst_s38417.g13175, inst_s38417.g12507, inst_s38417.g13182, inst_s38417.g13143, inst_s38417.g12524, inst_s38417.g13194, inst_s38417.g12457, inst_s38417.g12539, inst_s38417.g12467, inst_s38417.g12482, inst_s38417.g12499, inst_s38417.g13110, inst_s38417.g18669, inst_s38417.g18678, inst_s38417.g18707, inst_s38417.g18719, inst_s38417.g18726, inst_s38417.g18743, inst_s38417.g18755, inst_s38417.g18763, inst_s38417.g18780, inst_s38417.g18782, inst_s38417.g18794, inst_s38417.g18821, inst_s38417.g18804, inst_s38417.g18820, inst_s38417.g18835, inst_s38417.g18852, inst_s38417.g18836, inst_s38417.g18975, inst_s38417.g18837, inst_s38417.g18866, inst_s38417.g18968, inst_s38417.g18883, inst_s38417.g18867, inst_s38417.g18868, inst_s38417.g18885, inst_s38417.g18754, inst_s38417.g18906, inst_s38417.g18907, inst_s38417.g18781, inst_s38417.g18803, inst_s38417.g18942, inst_s38417.g18957, inst_s38417.g16654, inst_s38417.g16671, inst_s38417.g16692, inst_s38417.g16718, inst_s38417.g16860, inst_s38417.g16866, inst_s38417.g16803, inst_s38417.g16824, inst_s38417.g16835, inst_s38417.g16844, inst_s38417.g16845, inst_s38417.g16851, inst_s38417.g16853, inst_s38417.g16854, inst_s38417.g16857, inst_s38417.g16861, inst_s38417.g16880, inst_s38417.g16802, inst_s38417.g16823, inst_s38417.g17222, inst_s38417.g17224, inst_s38417.g17225, inst_s38417.g17226, inst_s38417.g17228, inst_s38417.g17229, inst_s38417.g17234, inst_s38417.g17235, inst_s38417.g17236, inst_s38417.g17246, inst_s38417.g17247, inst_s38417.g17248, inst_s38417.g17269, inst_s38417.g17270, inst_s38417.g17271, inst_s38417.g17302, inst_s38417.g17303, inst_s38417.g17340, inst_s38417.g17341, inst_s38417.g17383, inst_s38417.g17429, inst_s38417.g20310, inst_s38417.g20314, inst_s38417.g20333, inst_s38417.g20343, inst_s38417.g20353, inst_s38417.g20375, inst_s38417.g20376, inst_s38417.g20417, inst_s38417.g19144, inst_s38417.g19149, inst_s38417.g19153, inst_s38417.g19154, inst_s38417.g19157, inst_s38417.g19162, inst_s38417.g19163, inst_s38417.g19167, inst_s38417.g19172, inst_s38417.g19173, inst_s38417.g19178, inst_s38417.g19184, inst_s38417.g21842, inst_s38417.g21843, inst_s38417.g21845, inst_s38417.g21847, inst_s38417.g21851, inst_s38417.g21878, inst_s38417.g21880, inst_s38417.g21882, inst_s38417.g20874, inst_s38417.g20875, inst_s38417.g20876, inst_s38417.g20879, inst_s38417.g20880, inst_s38417.g20881, inst_s38417.g20882, inst_s38417.g20883, inst_s38417.g20682, inst_s38417.g20891, inst_s38417.g20892, inst_s38417.g20893, inst_s38417.g20894, inst_s38417.g20896, inst_s38417.g20897, inst_s38417.g20898, inst_s38417.g20899, inst_s38417.g20900, inst_s38417.g20901, inst_s38417.g20902, inst_s38417.g20903, inst_s38417.g20717, inst_s38417.g20910, inst_s38417.g20911, inst_s38417.g20912, inst_s38417.g20913, inst_s38417.g20915, inst_s38417.g20916, inst_s38417.g20917, inst_s38417.g20918, inst_s38417.g20919, inst_s38417.g20921, inst_s38417.g20922, inst_s38417.g20923, inst_s38417.g20924, inst_s38417.g20925, inst_s38417.g20926, inst_s38417.g20927, inst_s38417.g20752, inst_s38417.g20934, inst_s38417.g20935, inst_s38417.g20936, inst_s38417.g20937, inst_s38417.g20939, inst_s38417.g20940, inst_s38417.g20941, inst_s38417.g20944, inst_s38417.g20945, inst_s38417.g20946, inst_s38417.g20947, inst_s38417.g20948, inst_s38417.g20949, inst_s38417.g20950, inst_s38417.g20951, inst_s38417.g20952, inst_s38417.g20953, inst_s38417.g20954, inst_s38417.g20955, inst_s38417.g20789, inst_s38417.g20962, inst_s38417.g20963, inst_s38417.g20964, inst_s38417.g20965, inst_s38417.g20966, inst_s38417.g20967, inst_s38417.g20968, inst_s38417.g20969, inst_s38417.g20970, inst_s38417.g20972, inst_s38417.g20973, inst_s38417.g20974, inst_s38417.g20975, inst_s38417.g20976, inst_s38417.g20977, inst_s38417.g20978, inst_s38417.g20979, inst_s38417.g20980, inst_s38417.g20981, inst_s38417.g20982, inst_s38417.g20983, inst_s38417.g20989, inst_s38417.g20990, inst_s38417.g20991, inst_s38417.g20992, inst_s38417.g20993, inst_s38417.g20994, inst_s38417.g20995, inst_s38417.g20996, inst_s38417.g20997, inst_s38417.g20999, inst_s38417.g21000, inst_s38417.g21001, inst_s38417.g21002, inst_s38417.g21003, inst_s38417.g21004, inst_s38417.g21005, inst_s38417.g21006, inst_s38417.g21007, inst_s38417.g21009, inst_s38417.g21010, inst_s38417.g21011, inst_s38417.g21015, inst_s38417.g21016, inst_s38417.g21017, inst_s38417.g21018, inst_s38417.g21019, inst_s38417.g21020, inst_s38417.g21021, inst_s38417.g21022, inst_s38417.g21023, inst_s38417.g21025, inst_s38417.g21026, inst_s38417.g21027, inst_s38417.g21028, inst_s38417.g21029, inst_s38417.g21031, inst_s38417.g21032, inst_s38417.g21033, inst_s38417.g21034, inst_s38417.g21035, inst_s38417.g21039, inst_s38417.g21040, inst_s38417.g21041, inst_s38417.g21042, inst_s38417.g21043, inst_s38417.g21044, inst_s38417.g21045, inst_s38417.g21046, inst_s38417.g21047, inst_s38417.g21051, inst_s38417.g21052, inst_s38417.g21053, inst_s38417.g21054, inst_s38417.g21055, inst_s38417.g21056, inst_s38417.g21060, inst_s38417.g21061, inst_s38417.g21062, inst_s38417.g21063, inst_s38417.g21070, inst_s38417.g21071, inst_s38417.g21072, inst_s38417.g21073, inst_s38417.g21074, inst_s38417.g21075, inst_s38417.g21080, inst_s38417.g21081, inst_s38417.g21082, inst_s38417.g21094, inst_s38417.g20877, inst_s38417.g20884, inst_s38417.g21346, inst_s38417.g23000, inst_s38417.g23117, inst_s38417.g23014, inst_s38417.g23126, inst_s38417.g23022, inst_s38417.g23030, inst_s38417.g23137, inst_s38417.g23039, inst_s38417.g23047, inst_s38417.g21970, inst_s38417.g23058, inst_s38417.g23067, inst_s38417.g23076, inst_s38417.g23081, inst_s38417.g23092, inst_s38417.g23093, inst_s38417.g23097, inst_s38417.g23110, inst_s38417.g23111, inst_s38417.g23114, inst_s38417.g23123, inst_s38417.g23124, inst_s38417.g23132, inst_s38417.g23133, inst_s38417.g22025, inst_s38417.g22027, inst_s38417.g22028, inst_s38417.g22029, inst_s38417.g22030, inst_s38417.g22031, inst_s38417.g22032, inst_s38417.g22033, inst_s38417.g22034, inst_s38417.g22035, inst_s38417.g22037, inst_s38417.g22038, inst_s38417.g22039, inst_s38417.g22040, inst_s38417.g22041, inst_s38417.g22042, inst_s38417.g22043, inst_s38417.g22044, inst_s38417.g22045, inst_s38417.g22047, inst_s38417.g22048, inst_s38417.g22049, inst_s38417.g23136, inst_s38417.g22054, inst_s38417.g22055, inst_s38417.g22056, inst_s38417.g22057, inst_s38417.g22058, inst_s38417.g22059, inst_s38417.g22060, inst_s38417.g22061, inst_s38417.g22063, inst_s38417.g22064, inst_s38417.g22065, inst_s38417.g22066, inst_s38417.g22067, inst_s38417.g22068, inst_s38417.g21969, inst_s38417.g22073, inst_s38417.g22074, inst_s38417.g22075, inst_s38417.g22076, inst_s38417.g22077, inst_s38417.g22078, inst_s38417.g22079, inst_s38417.g22080, inst_s38417.g22081, inst_s38417.g22087, inst_s38417.g22088, inst_s38417.g22089, inst_s38417.g22090, inst_s38417.g22091, inst_s38417.g22092, inst_s38417.g21972, inst_s38417.g22097, inst_s38417.g22098, inst_s38417.g22099, inst_s38417.g22100, inst_s38417.g22101, inst_s38417.g22102, inst_s38417.g22103, inst_s38417.g22104, inst_s38417.g22105, inst_s38417.g22106, inst_s38417.g22112, inst_s38417.g22113, inst_s38417.g22114, inst_s38417.g22115, inst_s38417.g22116, inst_s38417.g22117, inst_s38417.g21974, inst_s38417.g22122, inst_s38417.g22123, inst_s38417.g22124, inst_s38417.g22125, inst_s38417.g22126, inst_s38417.g22127, inst_s38417.g22128, inst_s38417.g22129, inst_s38417.g22130, inst_s38417.g22131, inst_s38417.g22132, inst_s38417.g22138, inst_s38417.g22139, inst_s38417.g22140, inst_s38417.g22141, inst_s38417.g22142, inst_s38417.g22143, inst_s38417.g22145, inst_s38417.g22146, inst_s38417.g22147, inst_s38417.g22148, inst_s38417.g22149, inst_s38417.g22150, inst_s38417.g22151, inst_s38417.g22152, inst_s38417.g22153, inst_s38417.g22154, inst_s38417.g22155, inst_s38417.g22161, inst_s38417.g22162, inst_s38417.g22163, inst_s38417.g22164, inst_s38417.g22166, inst_s38417.g22167, inst_s38417.g22168, inst_s38417.g22169, inst_s38417.g22170, inst_s38417.g22171, inst_s38417.g22172, inst_s38417.g22173, inst_s38417.g22177, inst_s38417.g22178, inst_s38417.g22179, inst_s38417.g22180, inst_s38417.g22182, inst_s38417.g22183, inst_s38417.g22184, inst_s38417.g22185, inst_s38417.g22191, inst_s38417.g22192, inst_s38417.g22193, inst_s38417.g22194, inst_s38417.g22200, inst_s38417.g22578, inst_s38417.g22615, inst_s38417.g22651, inst_s38417.g22026, inst_s38417.g22218, inst_s38417.g22687, inst_s38417.g22231, inst_s38417.g22234, inst_s38417.g22242, inst_s38417.g22247, inst_s38417.g22249, inst_s38417.g22263, inst_s38417.g22267, inst_s38417.g22269, inst_s38417.g22280, inst_s38417.g22284, inst_s38417.g22299, inst_s38417.g23399, inst_s38417.g23406, inst_s38417.g24174, inst_s38417.g23413, inst_s38417.g24178, inst_s38417.g24179, inst_s38417.g23418, inst_s38417.g24181, inst_s38417.g24182, inst_s38417.g24206, inst_s38417.g24207, inst_s38417.g24208, inst_s38417.g24209, inst_s38417.g24212, inst_s38417.g24213, inst_s38417.g24214, inst_s38417.g24215, inst_s38417.g24216, inst_s38417.g24218, inst_s38417.g24219, inst_s38417.g24222, inst_s38417.g24223, inst_s38417.g24225, inst_s38417.g24226, inst_s38417.g24228, inst_s38417.g24230, inst_s38417.g24231, inst_s38417.g24235, inst_s38417.g24237, inst_s38417.g24238, inst_s38417.g24243, inst_s38417.g24250, inst_s38417.g23385, inst_s38417.g23392, inst_s38417.g23400, inst_s38417.g23324, inst_s38417.g23407, inst_s38417.g23329, inst_s38417.g23330, inst_s38417.g23339, inst_s38417.g23348, inst_s38417.g23357, inst_s38417.g23358, inst_s38417.g23359, inst_s38417.g24059, inst_s38417.g24072, inst_s38417.g24083, inst_s38417.g24092, inst_s38417.g25027, inst_s38417.g25042, inst_s38417.g25056, inst_s38417.g25067, inst_s38417.g24426, inst_s38417.g24430, inst_s38417.g24434, inst_s38417.g24438, inst_s38417.g24491, inst_s38417.g24498, inst_s38417.g24499, inst_s38417.g24501, inst_s38417.g24507, inst_s38417.g24508, inst_s38417.g24510, inst_s38417.g24511, inst_s38417.g24513, inst_s38417.g24445, inst_s38417.g24446, inst_s38417.g24519, inst_s38417.g24521, inst_s38417.g24522, inst_s38417.g24524, inst_s38417.g24525, inst_s38417.g24527, inst_s38417.g24532, inst_s38417.g24534, inst_s38417.g24535, inst_s38417.g24537, inst_s38417.g24538, inst_s38417.g24545, inst_s38417.g24547, inst_s38417.g24548, inst_s38417.g24557, inst_s38417.g24473, inst_s38417.g24476, inst_s38417.g25932, inst_s38417.g25935, inst_s38417.g25938, inst_s38417.g25940, inst_s38417.g25204, inst_s38417.g25206, inst_s38417.g25207, inst_s38417.g25209, inst_s38417.g25211, inst_s38417.g25212, inst_s38417.g25213, inst_s38417.g25214, inst_s38417.g25215, inst_s38417.g25217, inst_s38417.g25218, inst_s38417.g25219, inst_s38417.g25220, inst_s38417.g25221, inst_s38417.g25222, inst_s38417.g25223, inst_s38417.g25224, inst_s38417.g25225, inst_s38417.g25227, inst_s38417.g25228, inst_s38417.g25229, inst_s38417.g25230, inst_s38417.g25231, inst_s38417.g25232, inst_s38417.g25233, inst_s38417.g25234, inst_s38417.g25235, inst_s38417.g25236, inst_s38417.g25237, inst_s38417.g25239, inst_s38417.g25240, inst_s38417.g25241, inst_s38417.g25242, inst_s38417.g25243, inst_s38417.g25244, inst_s38417.g25245, inst_s38417.g25246, inst_s38417.g25247, inst_s38417.g25248, inst_s38417.g25249, inst_s38417.g25250, inst_s38417.g25251, inst_s38417.g25252, inst_s38417.g25253, inst_s38417.g25185, inst_s38417.g25255, inst_s38417.g25256, inst_s38417.g25257, inst_s38417.g25189, inst_s38417.g25259, inst_s38417.g25265, inst_s38417.g25191, inst_s38417.g25260, inst_s38417.g25194, inst_s38417.g25262, inst_s38417.g25263, inst_s38417.g25197, inst_s38417.g25266, inst_s38417.g25267, inst_s38417.g25268, inst_s38417.g25270, inst_s38417.g25271, inst_s38417.g25272, inst_s38417.g25279, inst_s38417.g25280, inst_s38417.g25199, inst_s38417.g25288, inst_s38417.g25201, inst_s38417.g25202, inst_s38417.g25450, inst_s38417.g25451, inst_s38417.g25452, inst_s38417.g26541, inst_s38417.g26545, inst_s38417.g26547, inst_s38417.g26553, inst_s38417.g26557, inst_s38417.g26559, inst_s38417.g26569, inst_s38417.g26573, inst_s38417.g26575, inst_s38417.g26592, inst_s38417.g26596, inst_s38417.g26616, inst_s38417.g26529, inst_s38417.g26530, inst_s38417.g26655, inst_s38417.g26531, inst_s38417.g26659, inst_s38417.g26661, inst_s38417.g26532, inst_s38417.g26664, inst_s38417.g26665, inst_s38417.g26667, inst_s38417.g26669, inst_s38417.g26670, inst_s38417.g26672, inst_s38417.g26675, inst_s38417.g26676, inst_s38417.g26025, inst_s38417.g26660, inst_s38417.g26666, inst_s38417.g26671, inst_s38417.g26677, inst_s38417.g26048, inst_s38417.g26031, inst_s38417.g26037, inst_s38417.g26183, inst_s38417.g27120, inst_s38417.g27123, inst_s38417.g27129, inst_s38417.g27131, inst_s38417.g26803, inst_s38417.g26804, inst_s38417.g26805, inst_s38417.g26806, inst_s38417.g26807, inst_s38417.g26808, inst_s38417.g26776, inst_s38417.g26809, inst_s38417.g26810, inst_s38417.g26811, inst_s38417.g26812, inst_s38417.g26813, inst_s38417.g26814, inst_s38417.g26781, inst_s38417.g26815, inst_s38417.g26816, inst_s38417.g26817, inst_s38417.g26786, inst_s38417.g26818, inst_s38417.g26820, inst_s38417.g26821, inst_s38417.g26789, inst_s38417.g26822, inst_s38417.g26823, inst_s38417.g26824, inst_s38417.g26825, inst_s38417.g26826, inst_s38417.g26795, inst_s38417.g26827, inst_s38417.g26798, inst_s38417.g27594, inst_s38417.g27603, inst_s38417.g27612, inst_s38417.g27621, inst_s38417.g27672, inst_s38417.g27678, inst_s38417.g27682, inst_s38417.g27243, inst_s38417.g27253, inst_s38417.g27255, inst_s38417.g27256, inst_s38417.g27257, inst_s38417.g27258, inst_s38417.g27259, inst_s38417.g27260, inst_s38417.g27261, inst_s38417.g27262, inst_s38417.g27263, inst_s38417.g27264, inst_s38417.g27265, inst_s38417.g27266, inst_s38417.g27267, inst_s38417.g27268, inst_s38417.g27269, inst_s38417.g27270, inst_s38417.g27271, inst_s38417.g27272, inst_s38417.g27273, inst_s38417.g27274, inst_s38417.g27275, inst_s38417.g27276, inst_s38417.g27277, inst_s38417.g27278, inst_s38417.g27279, inst_s38417.g27280, inst_s38417.g27281, inst_s38417.g27282, inst_s38417.g27283, inst_s38417.g27284, inst_s38417.g27285, inst_s38417.g27286, inst_s38417.g27287, inst_s38417.g27288, inst_s38417.g27289, inst_s38417.g27290, inst_s38417.g27291, inst_s38417.g27292, inst_s38417.g27293, inst_s38417.g27294, inst_s38417.g27295, inst_s38417.g27296, inst_s38417.g27297, inst_s38417.g27298, inst_s38417.g27299, inst_s38417.g27300, inst_s38417.g27301, inst_s38417.g27302, inst_s38417.g27303, inst_s38417.g27304, inst_s38417.g27305, inst_s38417.g27306, inst_s38417.g27307, inst_s38417.g27308, inst_s38417.g27309, inst_s38417.g27310, inst_s38417.g27311, inst_s38417.g27312, inst_s38417.g27313, inst_s38417.g27314, inst_s38417.g27315, inst_s38417.g27316, inst_s38417.g27317, inst_s38417.g27318, inst_s38417.g27319, inst_s38417.g27320, inst_s38417.g27321, inst_s38417.g27322, inst_s38417.g27323, inst_s38417.g27324, inst_s38417.g27325, inst_s38417.g27326, inst_s38417.g27327, inst_s38417.g27328, inst_s38417.g27329, inst_s38417.g27330, inst_s38417.g27331, inst_s38417.g27332, inst_s38417.g27333, inst_s38417.g27334, inst_s38417.g27335, inst_s38417.g27336, inst_s38417.g27337, inst_s38417.g27338, inst_s38417.g27339, inst_s38417.g27340, inst_s38417.g27341, inst_s38417.g27342, inst_s38417.g27343, inst_s38417.g27344, inst_s38417.g27345, inst_s38417.g27346, inst_s38417.g27347, inst_s38417.g27348, inst_s38417.g27354, inst_s38417.g28145, inst_s38417.g28146, inst_s38417.g28147, inst_s38417.g28148, inst_s38417.g28199, inst_s38417.g27718, inst_s38417.g27722, inst_s38417.g27724, inst_s38417.g27759, inst_s38417.g27760, inst_s38417.g27761, inst_s38417.g27762, inst_s38417.g27763, inst_s38417.g27764, inst_s38417.g27765, inst_s38417.g27766, inst_s38417.g27767, inst_s38417.g27768, inst_s38417.g27769, inst_s38417.g27771, inst_s38417.g28634, inst_s38417.g28635, inst_s38417.g28636, inst_s38417.g28637, inst_s38417.g28668, inst_s38417.g28321, inst_s38417.g28325, inst_s38417.g28328, inst_s38417.g28342, inst_s38417.g28344, inst_s38417.g28345, inst_s38417.g28346, inst_s38417.g28348, inst_s38417.g28349, inst_s38417.g28350, inst_s38417.g28351, inst_s38417.g28352, inst_s38417.g28353, inst_s38417.g28354, inst_s38417.g28355, inst_s38417.g28356, inst_s38417.g28357, inst_s38417.g28358, inst_s38417.g28360, inst_s38417.g28361, inst_s38417.g28362, inst_s38417.g28363, inst_s38417.g28364, inst_s38417.g28366, inst_s38417.g28367, inst_s38417.g28368, inst_s38417.g28371, inst_s38417.g28420, inst_s38417.g28421, inst_s38417.g28425, inst_s38417.g29109, inst_s38417.g29110, inst_s38417.g29111, inst_s38417.g29112, inst_s38417.g28732, inst_s38417.g28735, inst_s38417.g28736, inst_s38417.g28738, inst_s38417.g28744, inst_s38417.g28745, inst_s38417.g28746, inst_s38417.g28747, inst_s38417.g28749, inst_s38417.g28754, inst_s38417.g28758, inst_s38417.g28759, inst_s38417.g28760, inst_s38417.g28761, inst_s38417.g28990, inst_s38417.g28763, inst_s38417.g28767, inst_s38417.g28771, inst_s38417.g28772, inst_s38417.g28773, inst_s38417.g28774, inst_s38417.g28778, inst_s38417.g28782, inst_s38417.g28783, inst_s38417.g28788, inst_s38417.g28903, inst_s38417.g29353, inst_s38417.g29354, inst_s38417.g29355, inst_s38417.g29357, inst_s38417.g29167, inst_s38417.g29169, inst_s38417.g29170, inst_s38417.g29172, inst_s38417.g29173, inst_s38417.g29178, inst_s38417.g29179, inst_s38417.g29181, inst_s38417.g29182, inst_s38417.g29184, inst_s38417.g29185, inst_s38417.g29187, inst_s38417.g29194, inst_s38417.g29197, inst_s38417.g29198, inst_s38417.g29201, inst_s38417.g29204, inst_s38417.g29205, inst_s38417.g29209, inst_s38417.g29212, inst_s38417.g29213, inst_s38417.g29218, inst_s38417.g29221, inst_s38417.g29226, inst_s38417.g29579, inst_s38417.g29606, inst_s38417.g29608, inst_s38417.g29580, inst_s38417.g29609, inst_s38417.g29611, inst_s38417.g29612, inst_s38417.g29581, inst_s38417.g29613, inst_s38417.g29616, inst_s38417.g29617, inst_s38417.g29582, inst_s38417.g29618, inst_s38417.g29620, inst_s38417.g29621, inst_s38417.g29623, inst_s38417.g29936, inst_s38417.g29939, inst_s38417.g29941, inst_s38417.g30055, inst_s38417.g30072, inst_s38417.g30061, inst_s38417.g30267, inst_s38417.g30268, inst_s38417.g30269, inst_s38417.g30270, inst_s38417.g30271, inst_s38417.g30272, inst_s38417.g30273, inst_s38417.g30274, inst_s38417.g30275, inst_s38417.g30276, inst_s38417.g30277, inst_s38417.g30278, inst_s38417.g30279, inst_s38417.g30280, inst_s38417.g30281, inst_s38417.g30282, inst_s38417.g30283, inst_s38417.g30284, inst_s38417.g30285, inst_s38417.g30286, inst_s38417.g30287, inst_s38417.g30288, inst_s38417.g30289, inst_s38417.g30290, inst_s38417.g30291, inst_s38417.g30292, inst_s38417.g30293, inst_s38417.g30294, inst_s38417.g30295, inst_s38417.g30296, inst_s38417.g30297, inst_s38417.g30298, inst_s38417.g30299, inst_s38417.g30300, inst_s38417.g30301, inst_s38417.g30302, inst_s38417.g30303, inst_s38417.g30304, inst_s38417.g30245, inst_s38417.g30246, inst_s38417.g30247, inst_s38417.g30248, inst_s38417.g30249, inst_s38417.g30250, inst_s38417.g30251, inst_s38417.g30252, inst_s38417.g30253, inst_s38417.g30254, inst_s38417.g30255, inst_s38417.g30256, inst_s38417.g30257, inst_s38417.g30258, inst_s38417.g30259, inst_s38417.g30260, inst_s38417.g30261, inst_s38417.g30262, inst_s38417.g30263, inst_s38417.g30264, inst_s38417.g30265, inst_s38417.g30266, inst_s38417.g30455, inst_s38417.g30468, inst_s38417.g30470, inst_s38417.g30482, inst_s38417.g30485, inst_s38417.g30487, inst_s38417.g30500, inst_s38417.g30503, inst_s38417.g30505, inst_s38417.g30338, inst_s38417.g30341, inst_s38417.g30356, inst_s38417.g30668, inst_s38417.g30669, inst_s38417.g30670, inst_s38417.g30671, inst_s38417.g30672, inst_s38417.g30673, inst_s38417.g30674, inst_s38417.g30675, inst_s38417.g30676, inst_s38417.g30677, inst_s38417.g30678, inst_s38417.g30679, inst_s38417.g30680, inst_s38417.g30681, inst_s38417.g30682, inst_s38417.g30683, inst_s38417.g30684, inst_s38417.g30686, inst_s38417.g30687, inst_s38417.g30688, inst_s38417.g30689, inst_s38417.g30690, inst_s38417.g30691, inst_s38417.g30692, inst_s38417.g30693, inst_s38417.g30694, inst_s38417.g30695, inst_s38417.g30699, inst_s38417.g30700, inst_s38417.g30701, inst_s38417.g30702, inst_s38417.g30703, inst_s38417.g30704, inst_s38417.g30705, inst_s38417.g30706, inst_s38417.g30707, inst_s38417.g30708, inst_s38417.g30709, inst_s38417.g30566, inst_s38417.g30635, inst_s38417.g30636, inst_s38417.g30637, inst_s38417.g30638, inst_s38417.g30639, inst_s38417.g30640, inst_s38417.g30641, inst_s38417.g30642, inst_s38417.g30643, inst_s38417.g30644, inst_s38417.g30645, inst_s38417.g30646, inst_s38417.g30647, inst_s38417.g30648, inst_s38417.g30649, inst_s38417.g30650, inst_s38417.g30651, inst_s38417.g30652, inst_s38417.g30653, inst_s38417.g30654, inst_s38417.g30655, inst_s38417.g30656, inst_s38417.g30657, inst_s38417.g30658, inst_s38417.g30659, inst_s38417.g30660, inst_s38417.g30661, inst_s38417.g30662, inst_s38417.g30663, inst_s38417.g30664, inst_s38417.g30665, inst_s38417.g30666, inst_s38417.g30667, inst_s38417.g30796, inst_s38417.g30798, inst_s38417.g30801, inst_s38417.DFF_1_n1, inst_s38417.DFF_2_n1, inst_s38417.DFF_15_n1, inst_s38417.DFF_16_n1, inst_s38417.DFF_18_n1, inst_s38417.DFF_131_n1, inst_s38417.DFF_132_n1, inst_s38417.DFF_134_n1, inst_s38417.DFF_140_n1, inst_s38417.DFF_142_n1, inst_s38417.DFF_144_n1, inst_s38417.DFF_146_n1, inst_s38417.DFF_149_n1, inst_s38417.DFF_155_n1, inst_s38417.DFF_156_n1, inst_s38417.DFF_299_n1, inst_s38417.DFF_301_n1, inst_s38417.DFF_303_n1, inst_s38417.DFF_305_n1, inst_s38417.DFF_307_n1, inst_s38417.DFF_309_n1, inst_s38417.DFF_311_n1, inst_s38417.DFF_313_n1, inst_s38417.DFF_328_n1, inst_s38417.DFF_444_n1, inst_s38417.DFF_445_n1, inst_s38417.DFF_446_n1, inst_s38417.DFF_447_n1, inst_s38417.DFF_448_n1, inst_s38417.DFF_449_n1, inst_s38417.DFF_453_n1, inst_s38417.DFF_649_n1, inst_s38417.DFF_651_n1, inst_s38417.DFF_653_n1, inst_s38417.DFF_655_n1, inst_s38417.DFF_657_n1, inst_s38417.DFF_659_n1, inst_s38417.DFF_661_n1, inst_s38417.DFF_663_n1, inst_s38417.DFF_783_n1, inst_s38417.DFF_792_n1, inst_s38417.DFF_794_n1, inst_s38417.DFF_795_n1, inst_s38417.DFF_796_n1, inst_s38417.DFF_797_n1, inst_s38417.DFF_798_n1, inst_s38417.DFF_799_n1, inst_s38417.DFF_803_n1, inst_s38417.DFF_999_n1, inst_s38417.DFF_1001_n1, inst_s38417.DFF_1003_n1, inst_s38417.DFF_1005_n1, inst_s38417.DFF_1007_n1, inst_s38417.DFF_1009_n1, inst_s38417.DFF_1011_n1, inst_s38417.DFF_1013_n1, inst_s38417.DFF_1099_n1, inst_s38417.DFF_1100_n1, inst_s38417.DFF_1133_n1, inst_s38417.DFF_1142_n1, inst_s38417.DFF_1144_n1, inst_s38417.DFF_1145_n1, inst_s38417.DFF_1146_n1, inst_s38417.DFF_1147_n1, inst_s38417.DFF_1148_n1, inst_s38417.DFF_1149_n1, inst_s38417.DFF_1153_n1, inst_s38417.DFF_1349_n1, inst_s38417.DFF_1351_n1, inst_s38417.DFF_1353_n1, inst_s38417.DFF_1355_n1, inst_s38417.DFF_1357_n1, inst_s38417.DFF_1359_n1, inst_s38417.DFF_1361_n1, inst_s38417.DFF_1363_n1, inst_s38417.DFF_1378_n1, inst_s38417.DFF_1449_n1, inst_s38417.DFF_1450_n1, inst_s38417.DFF_1494_n1, inst_s38417.DFF_1495_n1, inst_s38417.DFF_1496_n1, inst_s38417.DFF_1497_n1, inst_s38417.DFF_1498_n1, inst_s38417.DFF_1499_n1, inst_s38417.DFF_1503_n1, inst_s38417.DFF_1561_n1, inst_s38417.DFF_1562_n1, inst_s38417.DFF_1612_n1, inst_s38417.DFF_1616_n1, inst_s38417.DFF_1617_n1, inst_s38417.DFF_1618_n1, inst_s38417.DFF_1625_n1, inst_s38417.DFF_1626_n1, inst_s38417.DFF_1628_n1, inst_s38417.n1565, inst_s38417.n1566, inst_s38417.n1567, inst_s38417.n1568, inst_s38417.n1569, inst_s38417.n1570, inst_s38417.n1572, inst_s38417.n1573, inst_s38417.n1574, inst_s38417.n1575, inst_s38417.n1576, inst_s38417.n1577, inst_s38417.n1578, inst_s38417.n1579, inst_s38417.n1580, inst_s38417.n1581, inst_s38417.n1582, inst_s38417.n1583, inst_s38417.n1584, inst_s38417.n1585, inst_s38417.n1586, inst_s38417.n1587, inst_s38417.n1590, inst_s38417.n1591, inst_s38417.n1592, inst_s38417.n1593, inst_s38417.n1594, inst_s38417.n1595, inst_s38417.n1596, inst_s38417.n1597, inst_s38417.n1598, inst_s38417.n1599, inst_s38417.n1600, inst_s38417.n1601, inst_s38417.n1603, inst_s38417.n1604, inst_s38417.n1605, inst_s38417.n1606, inst_s38417.n1607, inst_s38417.n1608, inst_s38417.n1609, inst_s38417.n1610, inst_s38417.n1611, inst_s38417.n1612, inst_s38417.n1613, inst_s38417.n1614, inst_s38417.n1615, inst_s38417.n1616, inst_s38417.n1617, inst_s38417.n1618, inst_s38417.n1619, inst_s38417.n1626, inst_s38417.n1628, inst_s38417.n1629, inst_s38417.n1630, inst_s38417.n1631, inst_s38417.n1632, inst_s38417.n1633, inst_s38417.n1634, inst_s38417.n1635, inst_s38417.n1636, inst_s38417.n1638, inst_s38417.n1640, inst_s38417.n1642, inst_s38417.n1645, inst_s38417.n1649, inst_s38417.n1650, inst_s38417.n1651, inst_s38417.n1652, inst_s38417.n1653, inst_s38417.n1654, inst_s38417.n1655, inst_s38417.n1657, inst_s38417.n1659, inst_s38417.n1661, inst_s38417.n1664, inst_s38417.n1668, inst_s38417.n1669, inst_s38417.n1670, inst_s38417.n1671, inst_s38417.n1672, inst_s38417.n1673, inst_s38417.n1674, inst_s38417.n1676, inst_s38417.n1678, inst_s38417.n1680, inst_s38417.n1683, inst_s38417.n1687, inst_s38417.n1688, inst_s38417.n1689, inst_s38417.n1690, inst_s38417.n1691, inst_s38417.n1692, inst_s38417.n1693, inst_s38417.n1695, inst_s38417.n1697, inst_s38417.n1699, inst_s38417.n1702, inst_s38417.n1745, inst_s38417.n1746, inst_s38417.n1747, inst_s38417.n1748, inst_s38417.n1759, inst_s38417.n1760, inst_s38417.n1761, inst_s38417.n1762, inst_s38417.n1763, inst_s38417.n1764, inst_s38417.n1765, inst_s38417.n1766, inst_s38417.n1768, inst_s38417.n1769, inst_s38417.n1770, inst_s38417.n1771, inst_s38417.n1772, inst_s38417.n1773, inst_s38417.n1774, inst_s38417.n1776, inst_s38417.n1778, inst_s38417.n1780, inst_s38417.n1781, inst_s38417.n1782, inst_s38417.n1783, inst_s38417.n1784, inst_s38417.n1785, inst_s38417.n1787, inst_s38417.n1788, inst_s38417.n1789, inst_s38417.n1790, inst_s38417.n1791, inst_s38417.n1792, inst_s38417.n1793, inst_s38417.n1794, inst_s38417.n1795, inst_s38417.n1796, inst_s38417.n1797, inst_s38417.n1798, inst_s38417.n1799, inst_s38417.n1801, inst_s38417.n1802, inst_s38417.n1808, inst_s38417.n1809, inst_s38417.n1810, inst_s38417.n1811, inst_s38417.n1812, inst_s38417.n1813, inst_s38417.n1814, inst_s38417.n1815, inst_s38417.n1816, inst_s38417.n1817, inst_s38417.n1818, inst_s38417.n1819, inst_s38417.n1820, inst_s38417.n1821, inst_s38417.n1822, inst_s38417.n1823, inst_s38417.n1824, inst_s38417.n1825, inst_s38417.n1826, inst_s38417.n1828, inst_s38417.n1829, inst_s38417.n1832, inst_s38417.n1833, inst_s38417.n1840, inst_s38417.n1841, inst_s38417.n1842, inst_s38417.n1843, inst_s38417.n1845, inst_s38417.n1846, inst_s38417.n1847, inst_s38417.n1848, inst_s38417.n1849, inst_s38417.n1850, inst_s38417.n1851, inst_s38417.n1852, inst_s38417.n1853, inst_s38417.n1854, inst_s38417.n1855, inst_s38417.n1857, inst_s38417.n1859, inst_s38417.n1860, inst_s38417.n1873, inst_s38417.n1874, inst_s38417.n1875, inst_s38417.n1876, inst_s38417.n1877, inst_s38417.n1878, inst_s38417.n1880, inst_s38417.n1882, inst_s38417.n1884, inst_s38417.n1885, inst_s38417.n1886, inst_s38417.n1887, inst_s38417.n1888, inst_s38417.n1889, inst_s38417.n1890, inst_s38417.n1891, inst_s38417.n1892, inst_s38417.n1893, inst_s38417.n1894, inst_s38417.n1895, inst_s38417.n1896, inst_s38417.n1897, inst_s38417.n1898, inst_s38417.n1899, inst_s38417.n1900, inst_s38417.n1901, inst_s38417.n1902, inst_s38417.n1903, inst_s38417.n1905, inst_s38417.n1906, inst_s38417.n1912, inst_s38417.n1913, inst_s38417.n1914, inst_s38417.n1915, inst_s38417.n1916, inst_s38417.n1917, inst_s38417.n1918, inst_s38417.n1919, inst_s38417.n1920, inst_s38417.n1921, inst_s38417.n1922, inst_s38417.n1923, inst_s38417.n1924, inst_s38417.n1925, inst_s38417.n1926, inst_s38417.n1927, inst_s38417.n1928, inst_s38417.n1932, inst_s38417.n1933, inst_s38417.n1941, inst_s38417.n1942, inst_s38417.n1943, inst_s38417.n1944, inst_s38417.n1946, inst_s38417.n1947, inst_s38417.n1948, inst_s38417.n1949, inst_s38417.n1950, inst_s38417.n1951, inst_s38417.n1952, inst_s38417.n1953, inst_s38417.n1954, inst_s38417.n1955, inst_s38417.n1956, inst_s38417.n1958, inst_s38417.n1960, inst_s38417.n1961, inst_s38417.n1974, inst_s38417.n1975, inst_s38417.n1976, inst_s38417.n1977, inst_s38417.n1978, inst_s38417.n1979, inst_s38417.n1980, inst_s38417.n1982, inst_s38417.n1984, inst_s38417.n1986, inst_s38417.n1987, inst_s38417.n1988, inst_s38417.n1989, inst_s38417.n1990, inst_s38417.n1993, inst_s38417.n1994, inst_s38417.n1995, inst_s38417.n1996, inst_s38417.n1997, inst_s38417.n1998, inst_s38417.n1999, inst_s38417.n2000, inst_s38417.n2001, inst_s38417.n2002, inst_s38417.n2003, inst_s38417.n2004, inst_s38417.n2005, inst_s38417.n2007, inst_s38417.n2008, inst_s38417.n2014, inst_s38417.n2015, inst_s38417.n2016, inst_s38417.n2017, inst_s38417.n2018, inst_s38417.n2019, inst_s38417.n2020, inst_s38417.n2021, inst_s38417.n2022, inst_s38417.n2023, inst_s38417.n2024, inst_s38417.n2025, inst_s38417.n2026, inst_s38417.n2027, inst_s38417.n2028, inst_s38417.n2029, inst_s38417.n2030, inst_s38417.n2034, inst_s38417.n2035, inst_s38417.n2043, inst_s38417.n2044, inst_s38417.n2045, inst_s38417.n2046, inst_s38417.n2048, inst_s38417.n2049, inst_s38417.n2050, inst_s38417.n2051, inst_s38417.n2052, inst_s38417.n2053, inst_s38417.n2054, inst_s38417.n2055, inst_s38417.n2056, inst_s38417.n2057, inst_s38417.n2058, inst_s38417.n2060, inst_s38417.n2062, inst_s38417.n2063, inst_s38417.n2076, inst_s38417.n2077, inst_s38417.n2078, inst_s38417.n2079, inst_s38417.n2080, inst_s38417.n2081, inst_s38417.n2082, inst_s38417.n2084, inst_s38417.n2086, inst_s38417.n2088, inst_s38417.n2089, inst_s38417.n2090, inst_s38417.n2091, inst_s38417.n2092, inst_s38417.n2095, inst_s38417.n2096, inst_s38417.n2097, inst_s38417.n2098, inst_s38417.n2099, inst_s38417.n2100, inst_s38417.n2101, inst_s38417.n2102, inst_s38417.n2103, inst_s38417.n2104, inst_s38417.n2105, inst_s38417.n2106, inst_s38417.n2107, inst_s38417.n2109, inst_s38417.n2110, inst_s38417.n2116, inst_s38417.n2117, inst_s38417.n2118, inst_s38417.n2119, inst_s38417.n2120, inst_s38417.n2121, inst_s38417.n2122, inst_s38417.n2123, inst_s38417.n2124, inst_s38417.n2125, inst_s38417.n2126, inst_s38417.n2127, inst_s38417.n2128, inst_s38417.n2129, inst_s38417.n2130, inst_s38417.n2131, inst_s38417.n2132, inst_s38417.n2136, inst_s38417.n2137, inst_s38417.n2145, inst_s38417.n2146, inst_s38417.n2147, inst_s38417.n2148, inst_s38417.n2150, inst_s38417.n2151, inst_s38417.n2152, inst_s38417.n2153, inst_s38417.n2154, inst_s38417.n2155, inst_s38417.n2156, inst_s38417.n2157, inst_s38417.n2158, inst_s38417.n2159, inst_s38417.n2160, inst_s38417.n2162, inst_s38417.n2164, inst_s38417.n2165, inst_s38417.n2180, inst_s38417.n2185, inst_s38417.n2186, inst_s38417.n2187, inst_s38417.n2188, inst_s38417.n2189, inst_s38417.n2190, inst_s38417.n2191, inst_s38417.n2192, inst_s38417.n2193, inst_s38417.n2195, inst_s38417.n2196, inst_s38417.n2197, inst_s38417.n2198, inst_s38417.n2199, inst_s38417.n2200, inst_s38417.n2201, inst_s38417.n2202, inst_s38417.n2203, inst_s38417.n2204, inst_s38417.n2205, inst_s38417.n2206, inst_s38417.n2207, inst_s38417.n2208, inst_s38417.n2209, inst_s38417.n2210, inst_s38417.n2211, inst_s38417.n2212, inst_s38417.n2213, inst_s38417.n2214, inst_s38417.n2215, inst_s38417.n2216, inst_s38417.n2217, inst_s38417.n2218, inst_s38417.n2219, inst_s38417.n2220, inst_s38417.n2221, inst_s38417.n2222, inst_s38417.n2223, inst_s38417.n2224, inst_s38417.n2225, inst_s38417.n2226, inst_s38417.n2227, inst_s38417.n2228, inst_s38417.n2229, inst_s38417.n2230, inst_s38417.n2231, inst_s38417.n2232, inst_s38417.n2233, inst_s38417.n2234, inst_s38417.n2235, inst_s38417.n2236, inst_s38417.n2237, inst_s38417.n2238, inst_s38417.n2239, inst_s38417.n2240, inst_s38417.n2241, inst_s38417.n2243, inst_s38417.n2244, inst_s38417.n2245, inst_s38417.n2246, inst_s38417.n2247, inst_s38417.n2248, inst_s38417.n2249, inst_s38417.n2250, inst_s38417.n2251, inst_s38417.n2252, inst_s38417.n2253, inst_s38417.n2254, inst_s38417.n2255, inst_s38417.n2256, inst_s38417.n2257, inst_s38417.n2258, inst_s38417.n2259, inst_s38417.n2260, inst_s38417.n2261, inst_s38417.n2262, inst_s38417.n2263, inst_s38417.n2264, inst_s38417.n2265, inst_s38417.n2267, inst_s38417.n2268, inst_s38417.n2269, inst_s38417.n2270, inst_s38417.n2271, inst_s38417.n2272, inst_s38417.n2273, inst_s38417.n2274, inst_s38417.n2275, inst_s38417.n2276, inst_s38417.n2277, inst_s38417.n2278, inst_s38417.n2279, inst_s38417.n2280, inst_s38417.n2281, inst_s38417.n2282, inst_s38417.n2283, inst_s38417.n2284, inst_s38417.n2285, inst_s38417.n2286, inst_s38417.n2287, inst_s38417.n2288, inst_s38417.n2289, inst_s38417.n2290, inst_s38417.n2291, inst_s38417.n2292, inst_s38417.n2293, inst_s38417.n2294, inst_s38417.n2295, inst_s38417.n2296, inst_s38417.n2297, inst_s38417.n2298, inst_s38417.n2299, inst_s38417.n2300, inst_s38417.n2301, inst_s38417.n2302, inst_s38417.n2303, inst_s38417.n2304, inst_s38417.n2305, inst_s38417.n2306, inst_s38417.n2307, inst_s38417.n2308, inst_s38417.n2309, inst_s38417.n2310, inst_s38417.n2311, inst_s38417.n2312, inst_s38417.n2313, inst_s38417.n2315, inst_s38417.n2316, inst_s38417.n2317, inst_s38417.n2318, inst_s38417.n2319, inst_s38417.n2320, inst_s38417.n2321, inst_s38417.n2322, inst_s38417.n2323, inst_s38417.n2324, inst_s38417.n2325, inst_s38417.n2326, inst_s38417.n2327, inst_s38417.n2328, inst_s38417.n2329, inst_s38417.n2330, inst_s38417.n2331, inst_s38417.n2332, inst_s38417.n2333, inst_s38417.n2334, inst_s38417.n2335, inst_s38417.n2336, inst_s38417.n2337, inst_s38417.n2339, inst_s38417.n2340, inst_s38417.n2341, inst_s38417.n2342, inst_s38417.n2343, inst_s38417.n2344, inst_s38417.n2345, inst_s38417.n2346, inst_s38417.n2347, inst_s38417.n2348, inst_s38417.n2349, inst_s38417.n2350, inst_s38417.n2351, inst_s38417.n2352, inst_s38417.n2353, inst_s38417.n2354, inst_s38417.n2355, inst_s38417.n2356, inst_s38417.n2357, inst_s38417.n2358, inst_s38417.n2359, inst_s38417.n2360, inst_s38417.n2361, inst_s38417.n2362, inst_s38417.n2363, inst_s38417.n2364, inst_s38417.n2365, inst_s38417.n2366, inst_s38417.n2367, inst_s38417.n2368, inst_s38417.n2369, inst_s38417.n2370, inst_s38417.n2371, inst_s38417.n2372, inst_s38417.n2373, inst_s38417.n2374, inst_s38417.n2375, inst_s38417.n2376, inst_s38417.n2377, inst_s38417.n2378, inst_s38417.n2379, inst_s38417.n2380, inst_s38417.n2381, inst_s38417.n2382, inst_s38417.n2383, inst_s38417.n2384, inst_s38417.n2385, inst_s38417.n2387, inst_s38417.n2388, inst_s38417.n2389, inst_s38417.n2390, inst_s38417.n2391, inst_s38417.n2392, inst_s38417.n2393, inst_s38417.n2394, inst_s38417.n2395, inst_s38417.n2396, inst_s38417.n2397, inst_s38417.n2398, inst_s38417.n2399, inst_s38417.n2400, inst_s38417.n2401, inst_s38417.n2402, inst_s38417.n2403, inst_s38417.n2404, inst_s38417.n2405, inst_s38417.n2406, inst_s38417.n2407, inst_s38417.n2408, inst_s38417.n2409, inst_s38417.n2410, inst_s38417.n2411, inst_s38417.n2412, inst_s38417.n2413, inst_s38417.n2414, inst_s38417.n2416, inst_s38417.n2417, inst_s38417.n2418, inst_s38417.n2419, inst_s38417.n2420, inst_s38417.n2421, inst_s38417.n2422, inst_s38417.n2423, inst_s38417.n2424, inst_s38417.n2425, inst_s38417.n2426, inst_s38417.n2427, inst_s38417.n2428, inst_s38417.n2429, inst_s38417.n2430, inst_s38417.n2431, inst_s38417.n2432, inst_s38417.n2433, inst_s38417.n2434, inst_s38417.n2435, inst_s38417.n2436, inst_s38417.n2437, inst_s38417.n2438, inst_s38417.n2439, inst_s38417.n2440, inst_s38417.n2441, inst_s38417.n2442, inst_s38417.n2443, inst_s38417.n2444, inst_s38417.n2445, inst_s38417.n2446, inst_s38417.n2447, inst_s38417.n2448, inst_s38417.n2450, inst_s38417.n2451, inst_s38417.n2452, inst_s38417.n2453, inst_s38417.n2454, inst_s38417.n2455, inst_s38417.n2456, inst_s38417.n2457, inst_s38417.n2458, inst_s38417.n2459, inst_s38417.n2460, inst_s38417.n2461, inst_s38417.n2462, inst_s38417.n2463, inst_s38417.n2464, inst_s38417.n2465, inst_s38417.n2466, inst_s38417.n2467, inst_s38417.n2468, inst_s38417.n2469, inst_s38417.n2470, inst_s38417.n2471, inst_s38417.n2472, inst_s38417.n2473, inst_s38417.n2474, inst_s38417.n2475, inst_s38417.n2476, inst_s38417.n2477, inst_s38417.n2478, inst_s38417.n2479, inst_s38417.n2480, inst_s38417.n2481, inst_s38417.n2482, inst_s38417.n2483, inst_s38417.n2484, inst_s38417.n2485, inst_s38417.n2486, inst_s38417.n2487, inst_s38417.n2488, inst_s38417.n2489, inst_s38417.n2490, inst_s38417.n2491, inst_s38417.n2492, inst_s38417.n2493, inst_s38417.n2494, inst_s38417.n2495, inst_s38417.n2496, inst_s38417.n2497, inst_s38417.n2498, inst_s38417.n2499, inst_s38417.n2500, inst_s38417.n2501, inst_s38417.n2502, inst_s38417.n2503, inst_s38417.n2504, inst_s38417.n2505, inst_s38417.n2506, inst_s38417.n2507, inst_s38417.n2508, inst_s38417.n2509, inst_s38417.n2510, inst_s38417.n2511, inst_s38417.n2512, inst_s38417.n2513, inst_s38417.n2514, inst_s38417.n2515, inst_s38417.n2516, inst_s38417.n2517, inst_s38417.n2518, inst_s38417.n2519, inst_s38417.n2520, inst_s38417.n2521, inst_s38417.n2522, inst_s38417.n2523, inst_s38417.n2524, inst_s38417.n2525, inst_s38417.n2526, inst_s38417.n2527, inst_s38417.n2528, inst_s38417.n2529, inst_s38417.n2530, inst_s38417.n2531, inst_s38417.n2532, inst_s38417.n2533, inst_s38417.n2534, inst_s38417.n2535, inst_s38417.n2536, inst_s38417.n2537, inst_s38417.n2538, inst_s38417.n2539, inst_s38417.n2540, inst_s38417.n2541, inst_s38417.n2542, inst_s38417.n2543, inst_s38417.n2544, inst_s38417.n2545, inst_s38417.n2546, inst_s38417.n2547, inst_s38417.n2548, inst_s38417.n2549, inst_s38417.n2550, inst_s38417.n2551, inst_s38417.n2552, inst_s38417.n2553, inst_s38417.n2554, inst_s38417.n2555, inst_s38417.n2556, inst_s38417.n2557, inst_s38417.n2558, inst_s38417.n2559, inst_s38417.n2560, inst_s38417.n2561, inst_s38417.n2562, inst_s38417.n2563, inst_s38417.n2564, inst_s38417.n2565, inst_s38417.n2566, inst_s38417.n2567, inst_s38417.n2568, inst_s38417.n2569, inst_s38417.n2570, inst_s38417.n2571, inst_s38417.n2572, inst_s38417.n2573, inst_s38417.n2574, inst_s38417.n2575, inst_s38417.n2576, inst_s38417.n2577, inst_s38417.n2578, inst_s38417.n2579, inst_s38417.n2580, inst_s38417.n2581, inst_s38417.n2582, inst_s38417.n2583, inst_s38417.n2584, inst_s38417.n2585, inst_s38417.n2586, inst_s38417.n2587, inst_s38417.n2588, inst_s38417.n2589, inst_s38417.n2590, inst_s38417.n2591, inst_s38417.n2592, inst_s38417.n2593, inst_s38417.n2594, inst_s38417.n2596, inst_s38417.n2597, inst_s38417.n2598, inst_s38417.n2599, inst_s38417.n2600, inst_s38417.n2601, inst_s38417.n2602, inst_s38417.n2603, inst_s38417.n2604, inst_s38417.n2605, inst_s38417.n2606, inst_s38417.n2607, inst_s38417.n2608, inst_s38417.n2609, inst_s38417.n2610, inst_s38417.n2611, inst_s38417.n2612, inst_s38417.n2613, inst_s38417.n2614, inst_s38417.n2615, inst_s38417.n2616, inst_s38417.n2617, inst_s38417.n2618, inst_s38417.n2619, inst_s38417.n2620, inst_s38417.n2621, inst_s38417.n2622, inst_s38417.n2623, inst_s38417.n2624, inst_s38417.n2625, inst_s38417.n2626, inst_s38417.n2627, inst_s38417.n2628, inst_s38417.n2629, inst_s38417.n2630, inst_s38417.n2631, inst_s38417.n2632, inst_s38417.n2633, inst_s38417.n2634, inst_s38417.n2635, inst_s38417.n2637, inst_s38417.n2638, inst_s38417.n2639, inst_s38417.n2640, inst_s38417.n2641, inst_s38417.n2642, inst_s38417.n2643, inst_s38417.n2644, inst_s38417.n2645, inst_s38417.n2646, inst_s38417.n2647, inst_s38417.n2648, inst_s38417.n2649, inst_s38417.n2650, inst_s38417.n2651, inst_s38417.n2652, inst_s38417.n2653, inst_s38417.n2654, inst_s38417.n2655, inst_s38417.n2656, inst_s38417.n2657, inst_s38417.n2658, inst_s38417.n2659, inst_s38417.n2660, inst_s38417.n2661, inst_s38417.n2662, inst_s38417.n2663, inst_s38417.n2664, inst_s38417.n2665, inst_s38417.n2666, inst_s38417.n2667, inst_s38417.n2668, inst_s38417.n2669, inst_s38417.n2670, inst_s38417.n2671, inst_s38417.n2672, inst_s38417.n2673, inst_s38417.n2674, inst_s38417.n2675, inst_s38417.n2676, inst_s38417.n2677, inst_s38417.n2678, inst_s38417.n2679, inst_s38417.n2680, inst_s38417.n2681, inst_s38417.n2682, inst_s38417.n2683, inst_s38417.n2684, inst_s38417.n2685, inst_s38417.n2686, inst_s38417.n2687, inst_s38417.n2688, inst_s38417.n2689, inst_s38417.n2690, inst_s38417.n2691, inst_s38417.n2692, inst_s38417.n2693, inst_s38417.n2694, inst_s38417.n2695, inst_s38417.n2696, inst_s38417.n2697, inst_s38417.n2698, inst_s38417.n2699, inst_s38417.n2700, inst_s38417.n2701, inst_s38417.n2702, inst_s38417.n2703, inst_s38417.n2704, inst_s38417.n2705, inst_s38417.n2706, inst_s38417.n2707, inst_s38417.n2708, inst_s38417.n2709, inst_s38417.n2710, inst_s38417.n2711, inst_s38417.n2712, inst_s38417.n2713, inst_s38417.n2714, inst_s38417.n2715, inst_s38417.n2716, inst_s38417.n2717, inst_s38417.n2718, inst_s38417.n2719, inst_s38417.n2720, inst_s38417.n2721, inst_s38417.n2722, inst_s38417.n2723, inst_s38417.n2724, inst_s38417.n2725, inst_s38417.n2726, inst_s38417.n2727, inst_s38417.n2728, inst_s38417.n2729, inst_s38417.n2730, inst_s38417.n2731, inst_s38417.n2732, inst_s38417.n2733, inst_s38417.n2734, inst_s38417.n2735, inst_s38417.n2736, inst_s38417.n2737, inst_s38417.n2738, inst_s38417.n2739, inst_s38417.n2740, inst_s38417.n2741, inst_s38417.n2742, inst_s38417.n2743, inst_s38417.n2744, inst_s38417.n2745, inst_s38417.n2746, inst_s38417.n2747, inst_s38417.n2748, inst_s38417.n2749, inst_s38417.n2750, inst_s38417.n2751, inst_s38417.n2752, inst_s38417.n2753, inst_s38417.n2754, inst_s38417.n2755, inst_s38417.n2756, inst_s38417.n2757, inst_s38417.n2758, inst_s38417.n2759, inst_s38417.n2760, inst_s38417.n2761, inst_s38417.n2762, inst_s38417.n2763, inst_s38417.n2764, inst_s38417.n2765, inst_s38417.n2766, inst_s38417.n2767, inst_s38417.n2768, inst_s38417.n2769, inst_s38417.n2770, inst_s38417.n2771, inst_s38417.n2772, inst_s38417.n2773, inst_s38417.n2774, inst_s38417.n2775, inst_s38417.n2777, inst_s38417.n2778, inst_s38417.n2779, inst_s38417.n2780, inst_s38417.n2781, inst_s38417.n2782, inst_s38417.n2783, inst_s38417.n2784, inst_s38417.n2785, inst_s38417.n2786, inst_s38417.n2787, inst_s38417.n2788, inst_s38417.n2789, inst_s38417.n2790, inst_s38417.n2791, inst_s38417.n2792, inst_s38417.n2793, inst_s38417.n2794, inst_s38417.n2795, inst_s38417.n2796, inst_s38417.n2797, inst_s38417.n2798, inst_s38417.n2799, inst_s38417.n2800, inst_s38417.n2801, inst_s38417.n2802, inst_s38417.n2803, inst_s38417.n2804, inst_s38417.n2805, inst_s38417.n2806, inst_s38417.n2807, inst_s38417.n2808, inst_s38417.n2809, inst_s38417.n2811, inst_s38417.n2812, inst_s38417.n2813, inst_s38417.n2814, inst_s38417.n2815, inst_s38417.n2816, inst_s38417.n2817, inst_s38417.n2818, inst_s38417.n2819, inst_s38417.n2821, inst_s38417.n2822, inst_s38417.n2823, inst_s38417.n2824, inst_s38417.n2825, inst_s38417.n2826, inst_s38417.n2827, inst_s38417.n2828, inst_s38417.n2829, inst_s38417.n2831, inst_s38417.n2832, inst_s38417.n2833, inst_s38417.n2834, inst_s38417.n2835, inst_s38417.n2836, inst_s38417.n2837, inst_s38417.n2838, inst_s38417.n2839, inst_s38417.n2840, inst_s38417.n2841, inst_s38417.n2842, inst_s38417.n2843, inst_s38417.n2844, inst_s38417.n2845, inst_s38417.n2846, inst_s38417.n2847, inst_s38417.n2848, inst_s38417.n2849, inst_s38417.n2850, inst_s38417.n2851, inst_s38417.n2852, inst_s38417.n2853, inst_s38417.n2854, inst_s38417.n2855, inst_s38417.n2856, inst_s38417.n2857, inst_s38417.n2858, inst_s38417.n2859, inst_s38417.n2860, inst_s38417.n2861, inst_s38417.n2862, inst_s38417.n2863, inst_s38417.n2864, inst_s38417.n2865, inst_s38417.n2866, inst_s38417.n2867, inst_s38417.n2868, inst_s38417.n2869, inst_s38417.n2870, inst_s38417.n2871, inst_s38417.n2872, inst_s38417.n2873, inst_s38417.n2874, inst_s38417.n2875, inst_s38417.n2876, inst_s38417.n2877, inst_s38417.n2878, inst_s38417.n2879, inst_s38417.n2880, inst_s38417.n2881, inst_s38417.n2882, inst_s38417.n2883, inst_s38417.n2884, inst_s38417.n2885, inst_s38417.n2886, inst_s38417.n2887, inst_s38417.n2888, inst_s38417.n2889, inst_s38417.n2890, inst_s38417.n2891, inst_s38417.n2892, inst_s38417.n2893, inst_s38417.n2894, inst_s38417.n2895, inst_s38417.n2896, inst_s38417.n2897, inst_s38417.n2898, inst_s38417.n2899, inst_s38417.n2900, inst_s38417.n2901, inst_s38417.n2902, inst_s38417.n2903, inst_s38417.n2904, inst_s38417.n2905, inst_s38417.n2906, inst_s38417.n2907, inst_s38417.n2908, inst_s38417.n2909, inst_s38417.n2910, inst_s38417.n2911, inst_s38417.n2912, inst_s38417.n2913, inst_s38417.n2914, inst_s38417.n2915, inst_s38417.n2916, inst_s38417.n2917, inst_s38417.n2918, inst_s38417.n2919, inst_s38417.n2920, inst_s38417.n2921, inst_s38417.n2922, inst_s38417.n2923, inst_s38417.n2924, inst_s38417.n2925, inst_s38417.n2926, inst_s38417.n2927, inst_s38417.n2928, inst_s38417.n2929, inst_s38417.n2930, inst_s38417.n2931, inst_s38417.n2932, inst_s38417.n2933, inst_s38417.n2934, inst_s38417.n2935, inst_s38417.n2936, inst_s38417.n2937, inst_s38417.n2938, inst_s38417.n2939, inst_s38417.n2940, inst_s38417.n2941, inst_s38417.n2942, inst_s38417.n2943, inst_s38417.n2944, inst_s38417.n2945, inst_s38417.n2946, inst_s38417.n2947, inst_s38417.n2948, inst_s38417.n2949, inst_s38417.n2950, inst_s38417.n2951, inst_s38417.n2952, inst_s38417.n2953, inst_s38417.n2954, inst_s38417.n2955, inst_s38417.n2956, inst_s38417.n2957, inst_s38417.n2958, inst_s38417.n2959, inst_s38417.n2960, inst_s38417.n2961, inst_s38417.n2963, inst_s38417.n2964, inst_s38417.n2965, inst_s38417.n2966, inst_s38417.n2967, inst_s38417.n2968, inst_s38417.n2969, inst_s38417.n2970, inst_s38417.n2971, inst_s38417.n2972, inst_s38417.n2973, inst_s38417.n2974, inst_s38417.n2975, inst_s38417.n2976, inst_s38417.n2977, inst_s38417.n2978, inst_s38417.n2979, inst_s38417.n2980, inst_s38417.n2981, inst_s38417.n2982, inst_s38417.n2983, inst_s38417.n2984, inst_s38417.n2985, inst_s38417.n2986, inst_s38417.n2987, inst_s38417.n2988, inst_s38417.n2989, inst_s38417.n2990, inst_s38417.n2991, inst_s38417.n2992, inst_s38417.n2993, inst_s38417.n2994, inst_s38417.n2995, inst_s38417.n2996, inst_s38417.n2997, inst_s38417.n2998, inst_s38417.n2999, inst_s38417.n3000, inst_s38417.n3001, inst_s38417.n3002, inst_s38417.n3003, inst_s38417.n3004, inst_s38417.n3005, inst_s38417.n3006, inst_s38417.n3007, inst_s38417.n3008, inst_s38417.n3009, inst_s38417.n3010, inst_s38417.n3011, inst_s38417.n3012, inst_s38417.n3013, inst_s38417.n3014, inst_s38417.n3015, inst_s38417.n3016, inst_s38417.n3017, inst_s38417.n3018, inst_s38417.n3019, inst_s38417.n3020, inst_s38417.n3021, inst_s38417.n3022, inst_s38417.n3023, inst_s38417.n3024, inst_s38417.n3025, inst_s38417.n3026, inst_s38417.n3027, inst_s38417.n3028, inst_s38417.n3029, inst_s38417.n3030, inst_s38417.n3031, inst_s38417.n3032, inst_s38417.n3033, inst_s38417.n3034, inst_s38417.n3035, inst_s38417.n3036, inst_s38417.n3037, inst_s38417.n3038, inst_s38417.n3039, inst_s38417.n3040, inst_s38417.n3041, inst_s38417.n3042, inst_s38417.n3043, inst_s38417.n3044, inst_s38417.n3045, inst_s38417.n3046, inst_s38417.n3047, inst_s38417.n3048, inst_s38417.n3049, inst_s38417.n3050, inst_s38417.n3051, inst_s38417.n3052, inst_s38417.n3053, inst_s38417.n3054, inst_s38417.n3055, inst_s38417.n3056, inst_s38417.n3057, inst_s38417.n3058, inst_s38417.n3059, inst_s38417.n3060, inst_s38417.n3061, inst_s38417.n3062, inst_s38417.n3063, inst_s38417.n3064, inst_s38417.n3065, inst_s38417.n3066, inst_s38417.n3067, inst_s38417.n3068, inst_s38417.n3069, inst_s38417.n3070, inst_s38417.n3071, inst_s38417.n3072, inst_s38417.n3073, inst_s38417.n3074, inst_s38417.n3075, inst_s38417.n3076, inst_s38417.n3077, inst_s38417.n3078, inst_s38417.n3079, inst_s38417.n3080, inst_s38417.n3081, inst_s38417.n3082, inst_s38417.n3083, inst_s38417.n3084, inst_s38417.n3085, inst_s38417.n3086, inst_s38417.n3087, inst_s38417.n3088, inst_s38417.n3089, inst_s38417.n3090, inst_s38417.n3091, inst_s38417.n3092, inst_s38417.n3093, inst_s38417.n3094, inst_s38417.n3095, inst_s38417.n3096, inst_s38417.n3097, inst_s38417.n3098, inst_s38417.n3099, inst_s38417.n3100, inst_s38417.n3101, inst_s38417.n3102, inst_s38417.n3103, inst_s38417.n3104, inst_s38417.n3105, inst_s38417.n3106, inst_s38417.n3107, inst_s38417.n3108, inst_s38417.n3109, inst_s38417.n3110, inst_s38417.n3111, inst_s38417.n3112, inst_s38417.n3113, inst_s38417.n3114, inst_s38417.n3115, inst_s38417.n3116, inst_s38417.n3117, inst_s38417.n3118, inst_s38417.n3119, inst_s38417.n3120, inst_s38417.n3121, inst_s38417.n3122, inst_s38417.n3123, inst_s38417.n3124, inst_s38417.n3125, inst_s38417.n3126, inst_s38417.n3127, inst_s38417.n3128, inst_s38417.n3129, inst_s38417.n3130, inst_s38417.n3131, inst_s38417.n3132, inst_s38417.n3133, inst_s38417.n3134, inst_s38417.n3135, inst_s38417.n3136, inst_s38417.n3137, inst_s38417.n3138, inst_s38417.n3139, inst_s38417.n3140, inst_s38417.n3141, inst_s38417.n3142, inst_s38417.n3143, inst_s38417.n3144, inst_s38417.n3145, inst_s38417.n3146, inst_s38417.n3147, inst_s38417.n3148, inst_s38417.n3149, inst_s38417.n3150, inst_s38417.n3151, inst_s38417.n3152, inst_s38417.n3153, inst_s38417.n3154, inst_s38417.n3155, inst_s38417.n3156, inst_s38417.n3157, inst_s38417.n3158, inst_s38417.n3159, inst_s38417.n3160, inst_s38417.n3161, inst_s38417.n3162, inst_s38417.n3163, inst_s38417.n3164, inst_s38417.n3165, inst_s38417.n3166, inst_s38417.n3167, inst_s38417.n3168, inst_s38417.n3169, inst_s38417.n3170, inst_s38417.n3171, inst_s38417.n3172, inst_s38417.n3173, inst_s38417.n3174, inst_s38417.n3176, inst_s38417.n3177, inst_s38417.n3178, inst_s38417.n3179, inst_s38417.n3180, inst_s38417.n3181, inst_s38417.n3182, inst_s38417.n3183, inst_s38417.n3184, inst_s38417.n3185, inst_s38417.n3186, inst_s38417.n3187, inst_s38417.n3188, inst_s38417.n3189, inst_s38417.n3190, inst_s38417.n3191, inst_s38417.n3192, inst_s38417.n3193, inst_s38417.n3194, inst_s38417.n3195, inst_s38417.n3196, inst_s38417.n3197, inst_s38417.n3198, inst_s38417.n3199, inst_s38417.n3200, inst_s38417.n3201, inst_s38417.n3202, inst_s38417.n3203, inst_s38417.n3204, inst_s38417.n3205, inst_s38417.n3206, inst_s38417.n3207, inst_s38417.n3208, inst_s38417.n3209, inst_s38417.n3210, inst_s38417.n3211, inst_s38417.n3212, inst_s38417.n3213, inst_s38417.n3214, inst_s38417.n3215, inst_s38417.n3216, inst_s38417.n3217, inst_s38417.n3218, inst_s38417.n3219, inst_s38417.n3220, inst_s38417.n3221, inst_s38417.n3222, inst_s38417.n3223, inst_s38417.n3224, inst_s38417.n3225, inst_s38417.n3226, inst_s38417.n3227, inst_s38417.n3228, inst_s38417.n3229, inst_s38417.n3230, inst_s38417.n3231, inst_s38417.n3232, inst_s38417.n3233, inst_s38417.n3234, inst_s38417.n3235, inst_s38417.n3236, inst_s38417.n3237, inst_s38417.n3238, inst_s38417.n3239, inst_s38417.n3240, inst_s38417.n3241, inst_s38417.n3242, inst_s38417.n3243, inst_s38417.n3244, inst_s38417.n3245, inst_s38417.n3246, inst_s38417.n3247, inst_s38417.n3248, inst_s38417.n3249, inst_s38417.n3250, inst_s38417.n3252, inst_s38417.n3253, inst_s38417.n3254, inst_s38417.n3255, inst_s38417.n3256, inst_s38417.n3257, inst_s38417.n3258, inst_s38417.n3259, inst_s38417.n3260, inst_s38417.n3261, inst_s38417.n3262, inst_s38417.n3263, inst_s38417.n3264, inst_s38417.n3265, inst_s38417.n3266, inst_s38417.n3267, inst_s38417.n3268, inst_s38417.n3269, inst_s38417.n3270, inst_s38417.n3271, inst_s38417.n3272, inst_s38417.n3273, inst_s38417.n3274, inst_s38417.n3275, inst_s38417.n3276, inst_s38417.n3277, inst_s38417.n3278, inst_s38417.n3279, inst_s38417.n3280, inst_s38417.n3281, inst_s38417.n3282, inst_s38417.n3283, inst_s38417.n3284, inst_s38417.n3285, inst_s38417.n3286, inst_s38417.n3287, inst_s38417.n3288, inst_s38417.n3289, inst_s38417.n3290, inst_s38417.n3291, inst_s38417.n3292, inst_s38417.n3293, inst_s38417.n3294, inst_s38417.n3295, inst_s38417.n3296, inst_s38417.n3297, inst_s38417.n3298, inst_s38417.n3299, inst_s38417.n3300, inst_s38417.n3301, inst_s38417.n3302, inst_s38417.n3303, inst_s38417.n3304, inst_s38417.n3305, inst_s38417.n3306, inst_s38417.n3307, inst_s38417.n3308, inst_s38417.n3309, inst_s38417.n3310, inst_s38417.n3311, inst_s38417.n3312, inst_s38417.n3313, inst_s38417.n3314, inst_s38417.n3315, inst_s38417.n3316, inst_s38417.n3317, inst_s38417.n3318, inst_s38417.n3319, inst_s38417.n3320, inst_s38417.n3321, inst_s38417.n3322, inst_s38417.n3323, inst_s38417.n3324, inst_s38417.n3325, inst_s38417.n3326, inst_s38417.n3327, inst_s38417.n3328, inst_s38417.n3329, inst_s38417.n3330, inst_s38417.n3331, inst_s38417.n3332, inst_s38417.n3333, inst_s38417.n3334, inst_s38417.n3335, inst_s38417.n3336, inst_s38417.n3337, inst_s38417.n3338, inst_s38417.n3339, inst_s38417.n3340, inst_s38417.n3341, inst_s38417.n3342, inst_s38417.n3343, inst_s38417.n3344, inst_s38417.n3345, inst_s38417.n3346, inst_s38417.n3347, inst_s38417.n3348, inst_s38417.n3349, inst_s38417.n3350, inst_s38417.n3351, inst_s38417.n3352, inst_s38417.n3353, inst_s38417.n3354, inst_s38417.n3355, inst_s38417.n3356, inst_s38417.n3357, inst_s38417.n3358, inst_s38417.n3359, inst_s38417.n3360, inst_s38417.n3361, inst_s38417.n3362, inst_s38417.n3363, inst_s38417.n3364, inst_s38417.n3365, inst_s38417.n3366, inst_s38417.n3367, inst_s38417.n3368, inst_s38417.n3369, inst_s38417.n3370, inst_s38417.n3371, inst_s38417.n3372, inst_s38417.n3373, inst_s38417.n3374, inst_s38417.n3375, inst_s38417.n3376, inst_s38417.n3377, inst_s38417.n3378, inst_s38417.n3379, inst_s38417.n3380, inst_s38417.n3381, inst_s38417.n3382, inst_s38417.n3383, inst_s38417.n3384, inst_s38417.n3385, inst_s38417.n3386, inst_s38417.n3387, inst_s38417.n3388, inst_s38417.n3389, inst_s38417.n3390, inst_s38417.n3391, inst_s38417.n3392, inst_s38417.n3393, inst_s38417.n3394, inst_s38417.n3395, inst_s38417.n3396, inst_s38417.n3397, inst_s38417.n3398, inst_s38417.n3399, inst_s38417.n3400, inst_s38417.n3401, inst_s38417.n3402, inst_s38417.n3403, inst_s38417.n3404, inst_s38417.n3405, inst_s38417.n3406, inst_s38417.n3407, inst_s38417.n3408, inst_s38417.n3409, inst_s38417.n3410, inst_s38417.n3411, inst_s38417.n3412, inst_s38417.n3413, inst_s38417.n3414, inst_s38417.n3415, inst_s38417.n3416, inst_s38417.n3417, inst_s38417.n3418, inst_s38417.n3419, inst_s38417.n3420, inst_s38417.n3421, inst_s38417.n3422, inst_s38417.n3423, inst_s38417.n3424, inst_s38417.n3425, inst_s38417.n3426, inst_s38417.n3427, inst_s38417.n3428, inst_s38417.n3429, inst_s38417.n3430, inst_s38417.n3431, inst_s38417.n3432, inst_s38417.n3433, inst_s38417.n3434, inst_s38417.n3435, inst_s38417.n3436, inst_s38417.n3437, inst_s38417.n3438, inst_s38417.n3439, inst_s38417.n3440, inst_s38417.n3441, inst_s38417.n3442, inst_s38417.n3443, inst_s38417.n3444, inst_s38417.n3445, inst_s38417.n3446, inst_s38417.n3447, inst_s38417.n3448, inst_s38417.n3449, inst_s38417.n3450, inst_s38417.n3451, inst_s38417.n3452, inst_s38417.n3453, inst_s38417.n3454, inst_s38417.n3455, inst_s38417.n3456, inst_s38417.n3457, inst_s38417.n3458, inst_s38417.n3459, inst_s38417.n3460, inst_s38417.n3461, inst_s38417.n3462, inst_s38417.n3463, inst_s38417.n3464, inst_s38417.n3465, inst_s38417.n3466, inst_s38417.n3467, inst_s38417.n3468, inst_s38417.n3469, inst_s38417.n3470, inst_s38417.n3471, inst_s38417.n3472, inst_s38417.n3473, inst_s38417.n3474, inst_s38417.n3475, inst_s38417.n3476, inst_s38417.n3477, inst_s38417.n3478, inst_s38417.n3479, inst_s38417.n3480, inst_s38417.n3481, inst_s38417.n3482, inst_s38417.n3483, inst_s38417.n3484, inst_s38417.n3485, inst_s38417.n3486, inst_s38417.n3487, inst_s38417.n3488, inst_s38417.n3489, inst_s38417.n3490, inst_s38417.n3491, inst_s38417.n3492, inst_s38417.n3493, inst_s38417.n3494, inst_s38417.n3495, inst_s38417.n3496, inst_s38417.n3497, inst_s38417.n3498, inst_s38417.n3499, inst_s38417.n3500, inst_s38417.n3501, inst_s38417.n3502, inst_s38417.n3503, inst_s38417.n3504, inst_s38417.n3505, inst_s38417.n3506, inst_s38417.n3507, inst_s38417.n3508, inst_s38417.n3509, inst_s38417.n3510, inst_s38417.n3511, inst_s38417.n3512, inst_s38417.n3513, inst_s38417.n3514, inst_s38417.n3515, inst_s38417.n3516, inst_s38417.n3517, inst_s38417.n3518, inst_s38417.n3519, inst_s38417.n3520, inst_s38417.n3521, inst_s38417.n3522, inst_s38417.n3523, inst_s38417.n3524, inst_s38417.n3525, inst_s38417.n3526, inst_s38417.n3527, inst_s38417.n3528, inst_s38417.n3529, inst_s38417.n3530, inst_s38417.n3531, inst_s38417.n3532, inst_s38417.n3533, inst_s38417.n3534, inst_s38417.n3535, inst_s38417.n3536, inst_s38417.n3537, inst_s38417.n3538, inst_s38417.n3539, inst_s38417.n3540, inst_s38417.n3541, inst_s38417.n3542, inst_s38417.n3543, inst_s38417.n3544, inst_s38417.n3545, inst_s38417.n3546, inst_s38417.n3547, inst_s38417.n3548, inst_s38417.n3549, inst_s38417.n3550, inst_s38417.n3551, inst_s38417.n3552, inst_s38417.n3553, inst_s38417.n3554, inst_s38417.n3555, inst_s38417.n3556, inst_s38417.n3557, inst_s38417.n3558, inst_s38417.n3559, inst_s38417.n3560, inst_s38417.n3561, inst_s38417.n3562, inst_s38417.n3563, inst_s38417.n3564, inst_s38417.n3565, inst_s38417.n3566, inst_s38417.n3567, inst_s38417.n3568, inst_s38417.n3569, inst_s38417.n3570, inst_s38417.n3571, inst_s38417.n3572, inst_s38417.n3573, inst_s38417.n3574, inst_s38417.n3575, inst_s38417.n3576, inst_s38417.n3577, inst_s38417.n3578, inst_s38417.n3579, inst_s38417.n3580, inst_s38417.n3581, inst_s38417.n3582, inst_s38417.n3583, inst_s38417.n3584, inst_s38417.n3585, inst_s38417.n3586, inst_s38417.n3587, inst_s38417.n3588, inst_s38417.n3589, inst_s38417.n3590, inst_s38417.n3591, inst_s38417.n3592, inst_s38417.n3593, inst_s38417.n3594, inst_s38417.n3595, inst_s38417.n3596, inst_s38417.n3597, inst_s38417.n3598, inst_s38417.n3599, inst_s38417.n3600, inst_s38417.n3601, inst_s38417.n3602, inst_s38417.n3603, inst_s38417.n3604, inst_s38417.n3605, inst_s38417.n3606, inst_s38417.n3607, inst_s38417.n3608, inst_s38417.n3609, inst_s38417.n3610, inst_s38417.n3611, inst_s38417.n3612, inst_s38417.n3613, inst_s38417.n3614, inst_s38417.n3615, inst_s38417.n3616, inst_s38417.n3617, inst_s38417.n3618, inst_s38417.n3619, inst_s38417.n3620, inst_s38417.n3621, inst_s38417.n3622, inst_s38417.n3623, inst_s38417.n3624, inst_s38417.n3625, inst_s38417.n3626, inst_s38417.n3627, inst_s38417.n3628, inst_s38417.n3629, inst_s38417.n3630, inst_s38417.n3631, inst_s38417.n3632, inst_s38417.n3633, inst_s38417.n3634, inst_s38417.n3635, inst_s38417.n3636, inst_s38417.n3637, inst_s38417.n3638, inst_s38417.n3639, inst_s38417.n3640, inst_s38417.n3641, inst_s38417.n3642, inst_s38417.n3643, inst_s38417.n3644, inst_s38417.n3645, inst_s38417.n3646, inst_s38417.n3647, inst_s38417.n3648, inst_s38417.n3649, inst_s38417.n3650, inst_s38417.n3651, inst_s38417.n3652, inst_s38417.n3653, inst_s38417.n3654, inst_s38417.n3655, inst_s38417.n3656, inst_s38417.n3657, inst_s38417.n3658, inst_s38417.n3659, inst_s38417.n3660, inst_s38417.n3661, inst_s38417.n3662, inst_s38417.n3663, inst_s38417.n3664, inst_s38417.n3665, inst_s38417.n3666, inst_s38417.n3667, inst_s38417.n3668, inst_s38417.n3669, inst_s38417.n3670, inst_s38417.n3671, inst_s38417.n3672, inst_s38417.n3673, inst_s38417.n3674, inst_s38417.n3675, inst_s38417.n3676, inst_s38417.n3677, inst_s38417.n3678, inst_s38417.n3679, inst_s38417.n3680, inst_s38417.n3681, inst_s38417.n3682, inst_s38417.n3683, inst_s38417.n3684, inst_s38417.n3685, inst_s38417.n3686, inst_s38417.n3687, inst_s38417.n3688, inst_s38417.n3689, inst_s38417.n3690, inst_s38417.n3691, inst_s38417.n3692, inst_s38417.n3693, inst_s38417.n3694, inst_s38417.n3695, inst_s38417.n3696, inst_s38417.n3697, inst_s38417.n3698, inst_s38417.n3699, inst_s38417.n3700, inst_s38417.n3701, inst_s38417.n3702, inst_s38417.n3703, inst_s38417.n3704, inst_s38417.n3705, inst_s38417.n3706, inst_s38417.n3707, inst_s38417.n3708, inst_s38417.n3709, inst_s38417.n3710, inst_s38417.n3711, inst_s38417.n3712, inst_s38417.n3713, inst_s38417.n3714, inst_s38417.n3715, inst_s38417.n3716, inst_s38417.n3718, inst_s38417.n3719, inst_s38417.n3720, inst_s38417.n3721, inst_s38417.n3722, inst_s38417.n3724, inst_s38417.n3725, inst_s38417.n3726, inst_s38417.n3727, inst_s38417.n3729, inst_s38417.n3730, inst_s38417.n3731, inst_s38417.n3733, inst_s38417.n3734, inst_s38417.n3735, inst_s38417.n3736, inst_s38417.n3737, inst_s38417.n3738, inst_s38417.n3739, inst_s38417.n3740, inst_s38417.n3741, inst_s38417.n3742, inst_s38417.n3743, inst_s38417.n3744, inst_s38417.n3745, inst_s38417.n3746, inst_s38417.n3747, inst_s38417.n3748, inst_s38417.n3749, inst_s38417.n3750, inst_s38417.n3751, inst_s38417.n3752, inst_s38417.n3753, inst_s38417.n3754, inst_s38417.n3755, inst_s38417.n3756, inst_s38417.n3757, inst_s38417.n3758, inst_s38417.n3759, inst_s38417.n3760, inst_s38417.n3761, inst_s38417.n3762, inst_s38417.n3763, inst_s38417.n3764, inst_s38417.n3765, inst_s38417.n3766, inst_s38417.n3767, inst_s38417.n3768, inst_s38417.n3769, inst_s38417.n3770, inst_s38417.n3771, inst_s38417.n3772, inst_s38417.n3773, inst_s38417.n3774, inst_s38417.n3775, inst_s38417.n3776, inst_s38417.n3777, inst_s38417.n3778, inst_s38417.n3781, inst_s38417.n3782, inst_s38417.n3783, inst_s38417.n3784, inst_s38417.n3785, inst_s38417.n3786, inst_s38417.n3787, inst_s38417.n3788, inst_s38417.n3789, inst_s38417.n3790, inst_s38417.n3791, inst_s38417.n3792, inst_s38417.n3793, inst_s38417.n3794, inst_s38417.n3795, inst_s38417.n3796, inst_s38417.n3797, inst_s38417.n3798, inst_s38417.n3799, inst_s38417.n3800, inst_s38417.n3801, inst_s38417.n3802, inst_s38417.n3803, inst_s38417.n3804, inst_s38417.n3805, inst_s38417.n3806, inst_s38417.n3807, inst_s38417.n3808, inst_s38417.n3811, inst_s38417.n3812, inst_s38417.n3813, inst_s38417.n3814, inst_s38417.n3815, inst_s38417.n3816, inst_s38417.n3817, inst_s38417.n3818, inst_s38417.n3819, inst_s38417.n3820, inst_s38417.n3821, inst_s38417.n3822, inst_s38417.n3823, inst_s38417.n3824, inst_s38417.n3825, inst_s38417.n3826, inst_s38417.n3827, inst_s38417.n3828, inst_s38417.n3829, inst_s38417.n3830, inst_s38417.n3831, inst_s38417.n3832, inst_s38417.n3833, inst_s38417.n3834, inst_s38417.n3835, inst_s38417.n3836, inst_s38417.n3839, inst_s38417.n3840, inst_s38417.n3841, inst_s38417.n3842, inst_s38417.n3843, inst_s38417.n3844, inst_s38417.n3845, inst_s38417.n3846, inst_s38417.n3847, inst_s38417.n3848, inst_s38417.n3850, inst_s38417.n3851, inst_s38417.n3852, inst_s38417.n3853, inst_s38417.n3854, inst_s38417.n3855, inst_s38417.n3857, inst_s38417.n3858, inst_s38417.n3859, inst_s38417.n3860, inst_s38417.n3861, inst_s38417.n3862, inst_s38417.n3863, inst_s38417.n3864, inst_s38417.n3865, inst_s38417.n3866, inst_s38417.n3867, inst_s38417.n3868, inst_s38417.n3869, inst_s38417.n3870, inst_s38417.n3871, inst_s38417.n3872, inst_s38417.n3873, inst_s38417.n3874, inst_s38417.n3875, inst_s38417.n3876, inst_s38417.n3877, inst_s38417.n3878, inst_s38417.n3879, inst_s38417.n3880, inst_s38417.n3881, inst_s38417.n3884, inst_s38417.n3885, inst_s38417.n3886, inst_s38417.n3887, inst_s38417.n3888, inst_s38417.n3889, inst_s38417.n3890, inst_s38417.n3891, inst_s38417.n3892, inst_s38417.n3893, inst_s38417.n3894, inst_s38417.n3895, inst_s38417.n3896, inst_s38417.n3897, inst_s38417.n3898, inst_s38417.n3899, inst_s38417.n3900, inst_s38417.n3901, inst_s38417.n3902, inst_s38417.n3903, inst_s38417.n3904, inst_s38417.n3905, inst_s38417.n3906, inst_s38417.n3907, inst_s38417.n3908, inst_s38417.n3909, inst_s38417.n3910, inst_s38417.n3911, inst_s38417.n3912, inst_s38417.n3913, inst_s38417.n3914, inst_s38417.n3915, inst_s38417.n3916, inst_s38417.n3917, inst_s38417.n3918, inst_s38417.n3919, inst_s38417.n3920, inst_s38417.n3921, inst_s38417.n3922, inst_s38417.n3923, inst_s38417.n3924, inst_s38417.n3925, inst_s38417.n3926, inst_s38417.n3927, inst_s38417.n3928, inst_s38417.n3929, inst_s38417.n3930, inst_s38417.n3931, inst_s38417.n3932, inst_s38417.n3933, inst_s38417.n3934, inst_s38417.n3935, inst_s38417.n3936, inst_s38417.n3937, inst_s38417.n3938, inst_s38417.n3939, inst_s38417.n3940, inst_s38417.n3941, inst_s38417.n3942, inst_s38417.n3943, inst_s38417.n3944, inst_s38417.n3945, inst_s38417.n3946, inst_s38417.n3947, inst_s38417.n3948, inst_s38417.n3949, inst_s38417.n3950, inst_s38417.n3951, inst_s38417.n3952, inst_s38417.n3953, inst_s38417.n3954, inst_s38417.n3955, inst_s38417.n3956, inst_s38417.n3957, inst_s38417.n3958, inst_s38417.n3959, inst_s38417.n3960, inst_s38417.n3961, inst_s38417.n3962, inst_s38417.n3963, inst_s38417.n3964, inst_s38417.n3965, inst_s38417.n3966, inst_s38417.n3967, inst_s38417.n3968, inst_s38417.n3969, inst_s38417.n3970, inst_s38417.n3971, inst_s38417.n3972, inst_s38417.n3973, inst_s38417.n3974, inst_s38417.n3975, inst_s38417.n3976, inst_s38417.n3977, inst_s38417.n3978, inst_s38417.n3979, inst_s38417.n3980, inst_s38417.n3981, inst_s38417.n3982, inst_s38417.n3983, inst_s38417.n3984, inst_s38417.n3985, inst_s38417.n3986, inst_s38417.n3987, inst_s38417.n3988, inst_s38417.n3989, inst_s38417.n3990, inst_s38417.n3991, inst_s38417.n3992, inst_s38417.n3993, inst_s38417.n3994, inst_s38417.n3995, inst_s38417.n3996, inst_s38417.n3997, inst_s38417.n3998, inst_s38417.n3999, inst_s38417.n4000, inst_s38417.n4001, inst_s38417.n4002, inst_s38417.n4003, inst_s38417.n4004, inst_s38417.n4005, inst_s38417.n4006, inst_s38417.n4007, inst_s38417.n4008, inst_s38417.n4009, inst_s38417.n4010, inst_s38417.n4011, inst_s38417.n4012, inst_s38417.n4013, inst_s38417.n4014, inst_s38417.n4015, inst_s38417.n4016, inst_s38417.n4017, inst_s38417.n4018, inst_s38417.n4019, inst_s38417.n4020, inst_s38417.n4021, inst_s38417.n4022, inst_s38417.n4023, inst_s38417.n4024, inst_s38417.n4025, inst_s38417.n4026, inst_s38417.n4027, inst_s38417.n4028, inst_s38417.n4029, inst_s38417.n4030, inst_s38417.n4031, inst_s38417.n4032, inst_s38417.n4033, inst_s38417.n4034, inst_s38417.n4035, inst_s38417.n4036, inst_s38417.n4037, inst_s38417.n4038, inst_s38417.n4039, inst_s38417.n4040, inst_s38417.n4041, inst_s38417.n4042, inst_s38417.n4043, inst_s38417.n4044, inst_s38417.n4045, inst_s38417.n4046, inst_s38417.n4047, inst_s38417.n4048, inst_s38417.n4049, inst_s38417.n4050, inst_s38417.n4051, inst_s38417.n4052, inst_s38417.n4053, inst_s38417.n4054, inst_s38417.n4055, inst_s38417.n4056, inst_s38417.n4057, inst_s38417.n4058, inst_s38417.n4059, inst_s38417.n4060, inst_s38417.n4061, inst_s38417.n4062, inst_s38417.n4063, inst_s38417.n4064, inst_s38417.n4065, inst_s38417.n4066, inst_s38417.n4067, inst_s38417.n4068, inst_s38417.n4069, inst_s38417.n4070, inst_s38417.n4071, inst_s38417.n4072, inst_s38417.n4073, inst_s38417.n4074, inst_s38417.n4075, inst_s38417.n4076, inst_s38417.n4077, inst_s38417.n4078, inst_s38417.n4079, inst_s38417.n4080, inst_s38417.n4081, inst_s38417.n4082, inst_s38417.n4083, inst_s38417.n4084, inst_s38417.n4085, inst_s38417.n4086, inst_s38417.n4087, inst_s38417.n4088, inst_s38417.n4089, inst_s38417.n4090, inst_s38417.n4091, inst_s38417.n4092, inst_s38417.n4093, inst_s38417.n4094, inst_s38417.n4095, inst_s38417.n4096, inst_s38417.n4097, inst_s38417.n4098, inst_s38417.n4099, inst_s38417.n4100, inst_s38417.n4101, inst_s38417.n4102, inst_s38417.n4103, inst_s38417.n4104, inst_s38417.n4105, inst_s38417.n4106, inst_s38417.n4107, inst_s38417.n4108, inst_s38417.n4109, inst_s38417.n4110, inst_s38417.n4111, inst_s38417.n4112, inst_s38417.n4113, inst_s38417.n4114, inst_s38417.n4115, inst_s38417.n4116, inst_s38417.n4117, inst_s38417.n4118, inst_s38417.n4119, inst_s38417.n4120, inst_s38417.n4121, inst_s38417.n4122, inst_s38417.n4123, inst_s38417.n4124, inst_s38417.n4125, inst_s38417.n4126, inst_s38417.n4127, inst_s38417.n4128, inst_s38417.n4129, inst_s38417.n4130, inst_s38417.n4131, inst_s38417.n4132, inst_s38417.n4133, inst_s38417.n4134, inst_s38417.n4135, inst_s38417.n4136, inst_s38417.n4137, inst_s38417.n4138, inst_s38417.n4139, inst_s38417.n4140, inst_s38417.n4141, inst_s38417.n4142, inst_s38417.n4143, inst_s38417.n4144, inst_s38417.n4145, inst_s38417.n4146, inst_s38417.n4147, inst_s38417.n4148, inst_s38417.n4149, inst_s38417.n4150, inst_s38417.n4151, inst_s38417.n4152, inst_s38417.n4153, inst_s38417.n4154, inst_s38417.n4155, inst_s38417.n4156, inst_s38417.n4157, inst_s38417.n4158, inst_s38417.n4159, inst_s38417.n4160, inst_s38417.n4161, inst_s38417.n4162, inst_s38417.n4163, inst_s38417.n4164, inst_s38417.n4165, inst_s38417.n4166, inst_s38417.n4167, inst_s38417.n4168, inst_s38417.n4169, inst_s38417.n4170, inst_s38417.n4171, inst_s38417.n4172, inst_s38417.n4173, inst_s38417.n4174, inst_s38417.n4175, inst_s38417.n4176, inst_s38417.n4177, inst_s38417.n4178, inst_s38417.n4179, inst_s38417.n4180, inst_s38417.n4181, inst_s38417.n4182, inst_s38417.n4183, inst_s38417.n4184, inst_s38417.n4185, inst_s38417.n4186, inst_s38417.n4187, inst_s38417.n4188, inst_s38417.n4189, inst_s38417.n4190, inst_s38417.n4191, inst_s38417.n4192, inst_s38417.n4193, inst_s38417.n4194, inst_s38417.n4195, inst_s38417.n4196, inst_s38417.n4197, inst_s38417.n4198, inst_s38417.n4199, inst_s38417.n4200, inst_s38417.n4201, inst_s38417.n4202, inst_s38417.n4203, inst_s38417.n4204, inst_s38417.n4205, inst_s38417.n4206, inst_s38417.n4207, inst_s38417.n4208, inst_s38417.n4210, inst_s38417.n4211, inst_s38417.n4212, inst_s38417.n4213, inst_s38417.n4214, inst_s38417.n4215, inst_s38417.n4216, inst_s38417.n4217, inst_s38417.n4218, inst_s38417.n4219, inst_s38417.n4220, inst_s38417.n4221, inst_s38417.n4222, inst_s38417.n4223, inst_s38417.n4224, inst_s38417.n4225, inst_s38417.n4226, inst_s38417.n4227, inst_s38417.n4228, inst_s38417.n4229, inst_s38417.n4230, inst_s38417.n4231, inst_s38417.n4232, inst_s38417.n4233, inst_s38417.n4234, inst_s38417.n4235, inst_s38417.n4236, inst_s38417.n4237, inst_s38417.n4238, inst_s38417.n4239, inst_s38417.n4240, inst_s38417.n4241, inst_s38417.n4242, inst_s38417.n4243, inst_s38417.n4244, inst_s38417.n4245, inst_s38417.n4246, inst_s38417.n4247, inst_s38417.n4248, inst_s38417.n4249, inst_s38417.n4250, inst_s38417.n4251, inst_s38417.n4252, inst_s38417.n4253, inst_s38417.n4254, inst_s38417.n4255, inst_s38417.n4256, inst_s38417.n4257, inst_s38417.n4258, inst_s38417.n4259, inst_s38417.n4260, inst_s38417.n4261, inst_s38417.n4262, inst_s38417.n4263, inst_s38417.n4264, inst_s38417.n4265, inst_s38417.n4266, inst_s38417.n4267, inst_s38417.n4268, inst_s38417.n4269, inst_s38417.n4270, inst_s38417.n4271, inst_s38417.n4272, inst_s38417.n4273, inst_s38417.n4274, inst_s38417.n4275, inst_s38417.n4276, inst_s38417.n4277, inst_s38417.n4278, inst_s38417.n4279, inst_s38417.n4280, inst_s38417.n4281, inst_s38417.n4282, inst_s38417.n4283, inst_s38417.n4284, inst_s38417.n4285, inst_s38417.n4287, inst_s38417.n4288, inst_s38417.n4289, inst_s38417.n4290, inst_s38417.n4291, inst_s38417.n4292, inst_s38417.n4293, inst_s38417.n4294, inst_s38417.n4295, inst_s38417.n4296, inst_s38417.n4297, inst_s38417.n4298, inst_s38417.n4299, inst_s38417.n4300, inst_s38417.n4301, inst_s38417.n4302, inst_s38417.n4303, inst_s38417.n4304, inst_s38417.n4305, inst_s38417.n4306, inst_s38417.n4307, inst_s38417.n4308, inst_s38417.n4309, inst_s38417.n4310, inst_s38417.n4311, inst_s38417.n4312, inst_s38417.n4313, inst_s38417.n4314, inst_s38417.n4315, inst_s38417.n4316, inst_s38417.n4317, inst_s38417.n4318, inst_s38417.n4319, inst_s38417.n4320, inst_s38417.n4321, inst_s38417.n4322, inst_s38417.n4323, inst_s38417.n4324, inst_s38417.n4325, inst_s38417.n4326, inst_s38417.n4327, inst_s38417.n4328, inst_s38417.n4329, inst_s38417.n4330, inst_s38417.n4331, inst_s38417.n4332, inst_s38417.n4333, inst_s38417.n4334, inst_s38417.n4335, inst_s38417.n4336, inst_s38417.n4337, inst_s38417.n4338, inst_s38417.n4339, inst_s38417.n4340, inst_s38417.n4341, inst_s38417.n4342, inst_s38417.n4343, inst_s38417.n4344, inst_s38417.n4345, inst_s38417.n4346, inst_s38417.n4347, inst_s38417.n4348, inst_s38417.n4349, inst_s38417.n4350, inst_s38417.n4351, inst_s38417.n4352, inst_s38417.n4353, inst_s38417.n4354, inst_s38417.n4355, inst_s38417.n4356, inst_s38417.n4357, inst_s38417.n4358, inst_s38417.n4359, inst_s38417.n4360, inst_s38417.n4361, inst_s38417.n4362, inst_s38417.n4363, inst_s38417.n4364, inst_s38417.n4365, inst_s38417.n4366, inst_s38417.n4367, inst_s38417.n4368, inst_s38417.n4369, inst_s38417.n4370, inst_s38417.n4371, inst_s38417.n4372, inst_s38417.n4373, inst_s38417.n4374, inst_s38417.n4375, inst_s38417.n4376, inst_s38417.n4377, inst_s38417.n4378, inst_s38417.n4379, inst_s38417.n4380, inst_s38417.n4381, inst_s38417.n4382, inst_s38417.n4383, inst_s38417.n4384, inst_s38417.n4385, inst_s38417.n4386, inst_s38417.n4387, inst_s38417.n4388, inst_s38417.n4389, inst_s38417.n4390, inst_s38417.n4391, inst_s38417.n4392, inst_s38417.n4393, inst_s38417.n4394, inst_s38417.n4395, inst_s38417.n4396, inst_s38417.n4397, inst_s38417.n4398, inst_s38417.n4399, inst_s38417.n4400, inst_s38417.n4401, inst_s38417.n4402, inst_s38417.n4403, inst_s38417.n4404, inst_s38417.n4405, inst_s38417.n4406, inst_s38417.n4407, inst_s38417.n4408, inst_s38417.n4409, inst_s38417.n4410, inst_s38417.n4411, inst_s38417.n4412, inst_s38417.n4413, inst_s38417.n4414, inst_s38417.n4415, inst_s38417.n4416, inst_s38417.n4417, inst_s38417.n4418, inst_s38417.n4419, inst_s38417.n4420, inst_s38417.n4421, inst_s38417.n4422, inst_s38417.n4423, inst_s38417.n4424, inst_s38417.n4425, inst_s38417.n4426, inst_s38417.n4427, inst_s38417.n4428, inst_s38417.n4429, inst_s38417.n4430, inst_s38417.n4431, inst_s38417.n4432, inst_s38417.n4433, inst_s38417.n4434, inst_s38417.n4435, inst_s38417.n4436, inst_s38417.n4437, inst_s38417.n4438, inst_s38417.n4439, inst_s38417.n4440, inst_s38417.n4441, inst_s38417.n4442, inst_s38417.n4443, inst_s38417.n4444, inst_s38417.n4445, inst_s38417.n4446, inst_s38417.n4447, inst_s38417.n4448, inst_s38417.n4449, inst_s38417.n4450, inst_s38417.n4451, inst_s38417.n4452, inst_s38417.n4453, inst_s38417.n4454, inst_s38417.n4455, inst_s38417.n4456, inst_s38417.n4457, inst_s38417.n4458, inst_s38417.n4459, inst_s38417.n4460, inst_s38417.n4461, inst_s38417.n4462, inst_s38417.n4463, inst_s38417.n4464, inst_s38417.n4465, inst_s38417.n4466, inst_s38417.n4467, inst_s38417.n4468, inst_s38417.n4469, inst_s38417.n4470, inst_s38417.n4471, inst_s38417.n4472, inst_s38417.n4473, inst_s38417.n4474, inst_s38417.n4475, inst_s38417.n4476, inst_s38417.n4477, inst_s38417.n4478, inst_s38417.n4479, inst_s38417.n4480, inst_s38417.n4481, inst_s38417.n4482, inst_s38417.n4483, inst_s38417.n4484, inst_s38417.n4485, inst_s38417.n4486, inst_s38417.n4487, inst_s38417.n4488, inst_s38417.n4489, inst_s38417.n4490, inst_s38417.n4491, inst_s38417.n4492, inst_s38417.n4493, inst_s38417.n4494, inst_s38417.n4495, inst_s38417.n4496, inst_s38417.n4497, inst_s38417.n4498, inst_s38417.n4499, inst_s38417.n4500, inst_s38417.n4501, inst_s38417.n4502, inst_s38417.n4503, inst_s38417.n4504, inst_s38417.n4505, inst_s38417.n4506, inst_s38417.n4507, inst_s38417.n4508, inst_s38417.n4509, inst_s38417.n4510, inst_s38417.n4511, inst_s38417.n4512, inst_s38417.n4513, inst_s38417.n4514, inst_s38417.n4515, inst_s38417.n4516, inst_s38417.n4517, inst_s38417.n4518, inst_s38417.n4519, inst_s38417.n4520, inst_s38417.n4521, inst_s38417.n4522, inst_s38417.n4523, inst_s38417.n4524, inst_s38417.n4525, inst_s38417.n4526, inst_s38417.n4527, inst_s38417.n4528, inst_s38417.n4529, inst_s38417.n4530, inst_s38417.n4531, inst_s38417.n4532, inst_s38417.n4533, inst_s38417.n4534, inst_s38417.n4535, inst_s38417.n4536, inst_s38417.n4537, inst_s38417.n4538, inst_s38417.n4539, inst_s38417.n4540, inst_s38417.n4541, inst_s38417.n4542, inst_s38417.n4543, inst_s38417.n4544, inst_s38417.n4545, inst_s38417.n4546, inst_s38417.n4547, inst_s38417.n4548, inst_s38417.n4549, inst_s38417.n4550, inst_s38417.n4551, inst_s38417.n4552, inst_s38417.n4553, inst_s38417.n4554, inst_s38417.n4555, inst_s38417.n4556, inst_s38417.n4557, inst_s38417.n4558, inst_s38417.n4559, inst_s38417.n4560, inst_s38417.n4561, inst_s38417.n4562, inst_s38417.n4563, inst_s38417.n4564, inst_s38417.n4565, inst_s38417.n4566, inst_s38417.n4567, inst_s38417.n4568, inst_s38417.n4569, inst_s38417.n4570, inst_s38417.n4571, inst_s38417.n4572, inst_s38417.n4573, inst_s38417.n4574, inst_s38417.n4575, inst_s38417.n4576, inst_s38417.n4577, inst_s38417.n4578, inst_s38417.n4579, inst_s38417.n4580, inst_s38417.n4581, inst_s38417.n4582, inst_s38417.n4583, inst_s38417.n4584, inst_s38417.n4585, inst_s38417.n4586, inst_s38417.n4587, inst_s38417.n4589, inst_s38417.n4591, inst_s38417.n4592, inst_s38417.n4593, inst_s38417.n4595, inst_s38417.n4596, inst_s38417.n4597, inst_s38417.n4598, inst_s38417.n4599, inst_s38417.n4600, inst_s38417.n4602, inst_s38417.n4604, inst_s38417.n4605, inst_s38417.n4606, inst_s38417.n4608, inst_s38417.n4610, inst_s38417.n4611, inst_s38417.n4612, inst_s38417.n4614, inst_s38417.n4616, inst_s38417.n4617, inst_s38417.n4618, inst_s38417.n4620, inst_s38417.n4622, inst_s38417.n4623, inst_s38417.n4624, inst_s38417.n4626, inst_s38417.n4628, inst_s38417.n4629, inst_s38417.n4630, inst_s38417.n4633, inst_s38417.n4634, inst_s38417.n4636, inst_s38417.n4638, inst_s38417.n4639, inst_s38417.n4640, inst_s38417.n4641, inst_s38417.n4643, inst_s38417.n4644, inst_s38417.n4646, inst_s38417.n4648, inst_s38417.n4649, inst_s38417.n4650, inst_s38417.n4651, inst_s38417.n4652, inst_s38417.n4653, inst_s38417.n4654, inst_s38417.n4655, inst_s38417.n4656, inst_s38417.n4657, inst_s38417.n4658, inst_s38417.n4659, inst_s38417.n4660, inst_s38417.n4661, inst_s38417.n4662, inst_s38417.n4663, inst_s38417.n4664, inst_s38417.n4665, inst_s38417.n4666, inst_s38417.n4667, inst_s38417.n4668, inst_s38417.n4669, inst_s38417.n4670, inst_s38417.n4671, inst_s38417.n4672, inst_s38417.n4673, inst_s38417.n4674, inst_s38417.n4675, inst_s38417.n4676, inst_s38417.n4677, inst_s38417.n4678, inst_s38417.n4679, inst_s38417.n4680, inst_s38417.n4681, inst_s38417.n4682, inst_s38417.n4683, inst_s38417.n4684, inst_s38417.n4685, inst_s38417.n4686, inst_s38417.n4687, inst_s38417.n4688, inst_s38417.n4689, inst_s38417.n4690, inst_s38417.n4691, inst_s38417.n4692, inst_s38417.n4693, inst_s38417.n4694, inst_s38417.n4695, inst_s38417.n4696, inst_s38417.n4697, inst_s38417.n4698, inst_s38417.n4699, inst_s38417.n4700, inst_s38417.n4701, inst_s38417.n4702, inst_s38417.n4703, inst_s38417.n4704, inst_s38417.n4705, inst_s38417.n4706, inst_s38417.n4707, inst_s38417.n4708, inst_s38417.n4709, inst_s38417.n4710, inst_s38417.n4711, inst_s38417.n4712, inst_s38417.n4713, inst_s38417.n4714, inst_s38417.n4715, inst_s38417.n4716, inst_s38417.n4717, inst_s38417.n4718, inst_s38417.n4719, inst_s38417.n4720, inst_s38417.n4721, inst_s38417.n4722, inst_s38417.n4723, inst_s38417.n4724, inst_s38417.n4725, inst_s38417.n4726, inst_s38417.n4727, inst_s38417.n4728, inst_s38417.n4729, inst_s38417.n4730, inst_s38417.n4731, inst_s38417.n4732, inst_s38417.n4733, inst_s38417.n4734, inst_s38417.n4735, inst_s38417.n4736, inst_s38417.n4737, inst_s38417.n4738, inst_s38417.n4739, inst_s38417.n4740, inst_s38417.n4741, inst_s38417.n4742, inst_s38417.n4743, inst_s38417.n4744, inst_s38417.n4745, inst_s38417.n4746, inst_s38417.n4747, inst_s38417.n4748, inst_s38417.n4749, inst_s38417.n4750, inst_s38417.n4751, inst_s38417.n4752, inst_s38417.n4753, inst_s38417.n4754, inst_s38417.n4755, inst_s38417.n4756, inst_s38417.n4757, inst_s38417.n4758, inst_s38417.n4759, inst_s38417.n4760, inst_s38417.n4761, inst_s38417.n4762, inst_s38417.n4763, inst_s38417.n4764, inst_s38417.n4765, inst_s38417.n4766, inst_s38417.n4767, inst_s38417.n4768, inst_s38417.n4769, inst_s38417.n4770, inst_s38417.n4771, inst_s38417.n4772, inst_s38417.n4773, inst_s38417.n4774, inst_s38417.n4775, inst_s38417.n4776, inst_s38417.n7907, inst_s38417.n7909, inst_s38417.n7912, inst_s38417.n7913, inst_s38417.n7918, inst_s38417.n7920, inst_s38417.n7921, inst_s38417.n7922, inst_s38417.n7923, inst_s38417.n7924, inst_s38417.n7925, inst_s38417.n7926, inst_s38417.n7929, inst_s38417.n7930, inst_s38417.n7936, inst_s38417.n7937, inst_s38417.n7938, inst_s38417.n7940, inst_s38417.n7941, inst_s38417.n7942, inst_s38417.n7943, inst_s38417.n7944, inst_s38417.n7945, inst_s38417.n7946, inst_s38417.n7960, inst_s38417.n7962, inst_s38417.n7963, inst_s38417.n7964, inst_s38417.n7965, inst_s38417.n7966, inst_s38417.n7967, inst_s38417.n7968, inst_s38417.n7971, inst_s38417.n7978, inst_s38417.n7979, inst_s38417.n7980, inst_s38417.n7983, inst_s38417.n7984, inst_s38417.n7985, inst_s38417.n7986, inst_s38417.n7987, inst_s38417.n7988, inst_s38417.n8003, inst_s38417.n8004, inst_s38417.n8005, inst_s38417.n8006, inst_s38417.n8007, inst_s38417.n8008, inst_s38417.n8009, inst_s38417.n8017, inst_s38417.n8018, inst_s38417.n8019, inst_s38417.n8020, inst_s38417.n8021, inst_s38417.n8024, inst_s38417.n8025, inst_s38417.n8026, inst_s38417.n8027, inst_s38417.n8040, inst_s38417.n8043, inst_s38417.n8044, inst_s38417.n8045, inst_s38417.n8046, inst_s38417.n8047, inst_s38417.n8055, inst_s38417.n8056, inst_s38417.n8057, inst_s38417.n8058, inst_s38417.n8059, inst_s38417.n8060, inst_s38417.n8061, inst_s38417.n8062, inst_s38417.n8065, inst_s38417.n8066, inst_s38417.n8076, inst_s38417.n8077, inst_s38417.n8078, inst_s38417.n8079, inst_s38417.n8080, inst_s38417.n8081, inst_s38417.n8082, inst_s38417.n8083, inst_s38417.n8084, inst_s38417.n8086, inst_s38417.n8087, inst_s38417.n8088, inst_s38417.n8089, inst_s38417.n8090, inst_s38417.n8098, inst_s38417.n8099, inst_s38417.n8102, inst_s38417.n8103, inst_s38417.n8104, inst_s38417.Tj_OUT1, inst_s38417.Tj_OUT1234, inst_s38417.Tj_OUT2, inst_s38417.Tj_OUT3, inst_s38417.Tj_OUT4, inst_s38417.Tj_OUT5, inst_s38417.Tj_OUT5678, inst_s38417.Tj_OUT6, inst_s38417.Tj_OUT7, inst_s38417.Tj_OUT8, inst_s38417.Tj_Payload, inst_s38417.Tj_Trigger, inst_s38417.n4263_Tj_Payload);
        end
        $fclose(fptr);
        $finish;
    end
endmodule